
module Cdf_Fetch ( clock, reset_n, start, ReadBus, ReadAddr, AccumlateOut, 
        StartOut, StoreAddress, input_base_offset, done );
  input [127:0] ReadBus;
  output [15:0] ReadAddr;
  output [19:0] AccumlateOut;
  output [15:0] StoreAddress;
  input clock, reset_n, start, input_base_offset;
  output StartOut, done;
  wire   n208, n210, \U3/U1/DATA1_1 , \U3/U1/DATA1_2 , \U3/U1/DATA1_3 ,
         \U3/U1/DATA1_4 , \U3/U1/DATA1_5 , \U3/U1/DATA1_6 , \U3/U1/DATA1_7 ,
         \U8/DATA1_0 , \U8/DATA1_1 , \U8/DATA1_2 , \U8/DATA1_3 , \U8/DATA1_4 ,
         \U8/DATA1_5 , \U8/DATA1_6 , \U8/DATA1_7 , \U8/DATA1_8 , \U8/DATA1_9 ,
         \U8/DATA1_10 , \U8/DATA1_11 , \U8/DATA1_12 , \U8/DATA1_13 ,
         \U8/DATA1_14 , \U8/DATA1_15 , \U8/DATA1_16 , \U8/DATA1_17 ,
         \U8/DATA1_18 , \U8/DATA1_19 , \U7/Z_0 , \U7/Z_1 , \U7/Z_2 , \U7/Z_3 ,
         \U7/Z_4 , \U7/Z_5 , \U7/Z_6 , \U7/Z_7 , \U7/Z_8 , \U7/Z_9 , \U7/Z_10 ,
         \U7/Z_11 , \U7/Z_12 , \U7/Z_13 , \U7/Z_14 , \U7/Z_15 , \U7/Z_16 ,
         \U7/Z_17 , \U7/Z_18 , \U7/Z_19 , \U5/Z_0 , \U5/Z_1 , \U5/Z_2 ,
         \U5/Z_3 , \U5/Z_4 , \U5/Z_5 , \U5/Z_6 , \U5/Z_7 , \U5/Z_8 , \U5/Z_9 ,
         \U5/Z_10 , \U5/Z_11 , \U5/Z_12 , \U5/Z_13 , \U5/Z_14 , \U4/Z_0 ,
         \U4/DATA3_0 , \add_63/carry[8] , \add_63/carry[7] , \add_63/carry[6] ,
         \add_63/carry[5] , \add_63/carry[4] , \add_63/carry[3] ,
         \add_63/carry[2] , \add_63/A[1] , \add_63/A[2] , \add_63/A[3] ,
         \add_63/A[4] , \add_63/A[5] , \add_63/A[6] , \add_63/A[7] ,
         \add_63/A[8] , \add_60/A[0] , \add_60/A[1] , \add_60/A[2] ,
         \add_60/A[3] , \add_60/A[4] , \add_60/A[5] , \add_60/A[6] ,
         \add_60/A[7] , \add_60/A[8] , \add_60/A[9] , \add_60/A[10] ,
         \add_60/A[11] , \add_60/A[12] , \add_60/A[13] , \add_60/A[14] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n36, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n375, n376,
         n377, n379, n381, n383, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n408, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446;
  assign \U8/DATA1_0  = ReadBus[0];
  assign \U8/DATA1_1  = ReadBus[1];
  assign \U8/DATA1_2  = ReadBus[2];
  assign \U8/DATA1_3  = ReadBus[3];
  assign \U8/DATA1_4  = ReadBus[4];
  assign \U8/DATA1_5  = ReadBus[5];
  assign \U8/DATA1_6  = ReadBus[6];
  assign \U8/DATA1_7  = ReadBus[7];
  assign \U8/DATA1_8  = ReadBus[8];
  assign \U8/DATA1_9  = ReadBus[9];
  assign \U8/DATA1_10  = ReadBus[10];
  assign \U8/DATA1_11  = ReadBus[11];
  assign \U8/DATA1_12  = ReadBus[12];
  assign \U8/DATA1_13  = ReadBus[13];
  assign \U8/DATA1_14  = ReadBus[14];
  assign \U8/DATA1_15  = ReadBus[15];
  assign \U8/DATA1_16  = ReadBus[16];
  assign \U8/DATA1_17  = ReadBus[17];
  assign \U8/DATA1_18  = ReadBus[18];
  assign \U8/DATA1_19  = ReadBus[19];
  assign \U4/DATA3_0  = input_base_offset;

  HA_X1 \add_63/U1_1_1  ( .A(\add_63/A[1] ), .B(n12), .CO(\add_63/carry[2] ), 
        .S(\U3/U1/DATA1_1 ) );
  HA_X1 \add_63/U1_1_2  ( .A(\add_63/A[2] ), .B(\add_63/carry[2] ), .CO(
        \add_63/carry[3] ), .S(\U3/U1/DATA1_2 ) );
  HA_X1 \add_63/U1_1_3  ( .A(\add_63/A[3] ), .B(\add_63/carry[3] ), .CO(
        \add_63/carry[4] ), .S(\U3/U1/DATA1_3 ) );
  HA_X1 \add_63/U1_1_4  ( .A(\add_63/A[4] ), .B(\add_63/carry[4] ), .CO(
        \add_63/carry[5] ), .S(\U3/U1/DATA1_4 ) );
  HA_X1 \add_63/U1_1_5  ( .A(\add_63/A[5] ), .B(\add_63/carry[5] ), .CO(
        \add_63/carry[6] ), .S(\U3/U1/DATA1_5 ) );
  HA_X1 \add_63/U1_1_6  ( .A(\add_63/A[6] ), .B(\add_63/carry[6] ), .CO(
        \add_63/carry[7] ), .S(\U3/U1/DATA1_6 ) );
  HA_X1 \add_63/U1_1_7  ( .A(\add_63/A[7] ), .B(\add_63/carry[7] ), .CO(
        \add_63/carry[8] ), .S(\U3/U1/DATA1_7 ) );
  TBUF_X2 \ReadAddr_tri[0]  ( .A(\add_60/A[0] ), .EN(n36), .Z(ReadAddr[0]) );
  TBUF_X2 \ReadAddr_tri[1]  ( .A(\add_60/A[1] ), .EN(n36), .Z(ReadAddr[1]) );
  TBUF_X2 \ReadAddr_tri[2]  ( .A(\add_60/A[2] ), .EN(n36), .Z(ReadAddr[2]) );
  TBUF_X2 \ReadAddr_tri[3]  ( .A(\add_60/A[3] ), .EN(n36), .Z(ReadAddr[3]) );
  TBUF_X2 \ReadAddr_tri[4]  ( .A(\add_60/A[4] ), .EN(n36), .Z(ReadAddr[4]) );
  TBUF_X2 \ReadAddr_tri[5]  ( .A(\add_60/A[5] ), .EN(n36), .Z(ReadAddr[5]) );
  TBUF_X2 \ReadAddr_tri[6]  ( .A(\add_60/A[6] ), .EN(n36), .Z(ReadAddr[6]) );
  TBUF_X2 \ReadAddr_tri[7]  ( .A(\add_60/A[7] ), .EN(n36), .Z(ReadAddr[7]) );
  TBUF_X2 \ReadAddr_tri[8]  ( .A(\add_60/A[8] ), .EN(n36), .Z(ReadAddr[8]) );
  TBUF_X2 \ReadAddr_tri[9]  ( .A(\add_60/A[9] ), .EN(n36), .Z(ReadAddr[9]) );
  TBUF_X2 \ReadAddr_tri[10]  ( .A(\add_60/A[10] ), .EN(n36), .Z(ReadAddr[10])
         );
  TBUF_X2 \ReadAddr_tri[11]  ( .A(\add_60/A[11] ), .EN(n36), .Z(ReadAddr[11])
         );
  TBUF_X2 \ReadAddr_tri[12]  ( .A(\add_60/A[12] ), .EN(n36), .Z(ReadAddr[12])
         );
  TBUF_X2 \ReadAddr_tri[13]  ( .A(\add_60/A[13] ), .EN(n36), .Z(ReadAddr[13])
         );
  TBUF_X2 \ReadAddr_tri[14]  ( .A(\add_60/A[14] ), .EN(n36), .Z(ReadAddr[14])
         );
  TBUF_X2 \ReadAddr_tri[15]  ( .A(n393), .EN(n36), .Z(ReadAddr[15]) );
  OAI22_X1 U3 ( .A1(n2), .A2(n3), .B1(n32), .B2(n4), .ZN(n40) );
  OAI22_X1 U5 ( .A1(n2), .A2(n5), .B1(n31), .B2(n4), .ZN(n41) );
  OAI22_X1 U7 ( .A1(n2), .A2(n6), .B1(n30), .B2(n4), .ZN(n42) );
  OAI22_X1 U9 ( .A1(n2), .A2(n7), .B1(n29), .B2(n4), .ZN(n43) );
  OAI22_X1 U11 ( .A1(n2), .A2(n8), .B1(n28), .B2(n4), .ZN(n44) );
  OAI22_X1 U13 ( .A1(n2), .A2(n9), .B1(n27), .B2(n4), .ZN(n45) );
  OAI22_X1 U15 ( .A1(n2), .A2(n10), .B1(n26), .B2(n4), .ZN(n46) );
  INV_X1 U18 ( .A(\add_63/carry[8] ), .ZN(n11) );
  OAI22_X1 U19 ( .A1(n2), .A2(n12), .B1(n47), .B2(n4), .ZN(n49) );
  AND2_X1 U30 ( .A1(\U8/DATA1_19 ), .A2(n375), .ZN(\U7/Z_19 ) );
  AND2_X1 U31 ( .A1(\U8/DATA1_18 ), .A2(n375), .ZN(\U7/Z_18 ) );
  AND2_X1 U32 ( .A1(\U8/DATA1_17 ), .A2(n375), .ZN(\U7/Z_17 ) );
  AND2_X1 U33 ( .A1(\U8/DATA1_16 ), .A2(n375), .ZN(\U7/Z_16 ) );
  AND2_X1 U34 ( .A1(\U8/DATA1_15 ), .A2(n375), .ZN(\U7/Z_15 ) );
  AND2_X1 U35 ( .A1(\U8/DATA1_14 ), .A2(n375), .ZN(\U7/Z_14 ) );
  NOR3_X1 U43 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n17) );
  NAND3_X1 U44 ( .A1(ReadBus[33]), .A2(ReadBus[31]), .A3(ReadBus[35]), .ZN(n20) );
  NAND3_X1 U45 ( .A1(ReadBus[27]), .A2(ReadBus[25]), .A3(ReadBus[29]), .ZN(n19) );
  NAND4_X1 U46 ( .A1(ReadBus[21]), .A2(start), .A3(ReadBus[23]), .A4(n21), 
        .ZN(n18) );
  NOR4_X1 U47 ( .A1(ReadBus[26]), .A2(ReadBus[24]), .A3(ReadBus[22]), .A4(
        ReadBus[20]), .ZN(n21) );
  NOR4_X1 U48 ( .A1(n22), .A2(ReadBus[39]), .A3(ReadBus[41]), .A4(ReadBus[40]), 
        .ZN(n16) );
  OR4_X1 U49 ( .A1(ReadBus[43]), .A2(ReadBus[42]), .A3(ReadBus[45]), .A4(
        ReadBus[44]), .ZN(n22) );
  NOR4_X1 U50 ( .A1(ReadBus[38]), .A2(ReadBus[37]), .A3(ReadBus[36]), .A4(
        ReadBus[34]), .ZN(n15) );
  NOR3_X1 U51 ( .A1(ReadBus[28]), .A2(ReadBus[32]), .A3(ReadBus[30]), .ZN(n14)
         );
  DFFR_X2 \AccumlateOut_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .RN(reset_n), .QN(
        n408) );
  DFFR_X2 \AccumlateOut_reg[0]  ( .D(\U7/Z_0 ), .CK(clock), .RN(reset_n), .QN(
        n406) );
  DFFR_X2 \AccumlateOut_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .RN(n414), .Q(
        AccumlateOut[2]) );
  DFFR_X2 \AccumlateOut_reg[5]  ( .D(\U7/Z_5 ), .CK(clock), .RN(n414), .QN(
        n381) );
  DFFR_X2 \AccumlateOut_reg[6]  ( .D(\U7/Z_6 ), .CK(clock), .RN(n414), .QN(
        n383) );
  DFFR_X2 \ReadAddress_reg[5]  ( .D(\U5/Z_5 ), .CK(clock), .RN(n411), .Q(
        \add_60/A[5] ), .QN(n399) );
  DFFR_X2 \ReadAddress_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .RN(n410), .Q(
        \add_60/A[2] ), .QN(n397) );
  DFFR_X2 \ReadAddress_reg[0]  ( .D(\U5/Z_0 ), .CK(clock), .RN(n410), .Q(
        \add_60/A[0] ), .QN(n33) );
  DFFR_X2 \ReadAddress_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .RN(n410), .Q(
        \add_60/A[1] ), .QN(n386) );
  DFFR_X2 \ReadAddress_reg[10]  ( .D(\U5/Z_10 ), .CK(clock), .RN(n411), .Q(
        \add_60/A[10] ), .QN(n402) );
  DFFR_X2 \AccumlateOut_reg[7]  ( .D(\U7/Z_7 ), .CK(clock), .RN(n414), .QN(
        n379) );
  DFFR_X2 done0_reg ( .D(n377), .CK(clock), .RN(reset_n), .Q(n210) );
  DFFR_X2 StartOut_reg ( .D(n376), .CK(clock), .RN(reset_n), .Q(StartOut) );
  DFFR_X2 \ReadAddress_reg[3]  ( .D(\U5/Z_3 ), .CK(clock), .RN(n410), .Q(
        \add_60/A[3] ), .QN(n398) );
  DFFR_X2 \ReadAddress_reg[7]  ( .D(\U5/Z_7 ), .CK(clock), .RN(n411), .Q(
        \add_60/A[7] ), .QN(n400) );
  DFFR_X2 \count_reg[0]  ( .D(n49), .CK(clock), .RN(n412), .Q(n12), .QN(n47)
         );
  DFFR_X2 \count_reg[2]  ( .D(n41), .CK(clock), .RN(n413), .Q(\add_63/A[2] ), 
        .QN(n31) );
  DFFR_X2 \count_reg[1]  ( .D(n40), .CK(clock), .RN(n412), .Q(\add_63/A[1] ), 
        .QN(n32) );
  DFFR_X2 \count_reg[3]  ( .D(n42), .CK(clock), .RN(n413), .Q(\add_63/A[3] ), 
        .QN(n30) );
  DFFR_X2 \ReadAddress_reg[9]  ( .D(\U5/Z_9 ), .CK(clock), .RN(n411), .Q(
        \add_60/A[9] ), .QN(n401) );
  DFFR_X2 \count_reg[4]  ( .D(n43), .CK(clock), .RN(n413), .Q(\add_63/A[4] ), 
        .QN(n29) );
  DFFR_X2 \count_reg[5]  ( .D(n44), .CK(clock), .RN(n413), .Q(\add_63/A[5] ), 
        .QN(n28) );
  DFFR_X2 \ReadAddress_reg[11]  ( .D(\U5/Z_11 ), .CK(clock), .RN(n412), .Q(
        \add_60/A[11] ), .QN(n403) );
  DFFR_X2 \ReadAddress_reg[13]  ( .D(\U5/Z_13 ), .CK(clock), .RN(n412), .Q(
        \add_60/A[13] ), .QN(n405) );
  DFFR_X2 \count_reg[6]  ( .D(n45), .CK(clock), .RN(n413), .Q(\add_63/A[6] ), 
        .QN(n27) );
  DFFR_X2 \count_reg[8]  ( .D(n48), .CK(clock), .RN(n410), .Q(\add_63/A[8] ), 
        .QN(n1) );
  DFFR_X2 \ReadAddress_reg[12]  ( .D(\U5/Z_12 ), .CK(clock), .RN(n412), .Q(
        \add_60/A[12] ), .QN(n404) );
  DFFR_X2 \count_reg[7]  ( .D(n46), .CK(clock), .RN(n413), .Q(\add_63/A[7] ), 
        .QN(n26) );
  DFFR_X2 \ReadAddress_reg[15]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n412), .Q(n393), .QN(n34) );
  DFFR_X2 \AccumlateOut_reg[8]  ( .D(\U7/Z_8 ), .CK(clock), .RN(reset_n), .Q(
        AccumlateOut[8]) );
  DFFR_X2 done_reg ( .D(n208), .CK(clock), .RN(n410), .Q(done) );
  DFFR_X2 \ReadAddress_reg[4]  ( .D(\U5/Z_4 ), .CK(clock), .RN(n410), .Q(
        \add_60/A[4] ) );
  DFFR_X2 done1_reg ( .D(n210), .CK(clock), .RN(reset_n), .Q(n208) );
  DFFR_X2 \StoreAddress_reg[15]  ( .D(n393), .CK(clock), .RN(n412), .Q(
        StoreAddress[15]) );
  DFFR_X2 \StoreAddress_reg[0]  ( .D(\add_60/A[0] ), .CK(clock), .RN(n410), 
        .Q(StoreAddress[0]) );
  DFFR_X2 \StoreAddress_reg[10]  ( .D(\add_60/A[10] ), .CK(clock), .RN(n411), 
        .Q(StoreAddress[10]) );
  DFFR_X2 \StoreAddress_reg[5]  ( .D(\add_60/A[5] ), .CK(clock), .RN(n411), 
        .Q(StoreAddress[5]) );
  DFFR_X2 \StoreAddress_reg[2]  ( .D(\add_60/A[2] ), .CK(clock), .RN(n410), 
        .Q(StoreAddress[2]) );
  DFFR_X2 \StoreAddress_reg[1]  ( .D(\add_60/A[1] ), .CK(clock), .RN(n410), 
        .Q(StoreAddress[1]) );
  DFFR_X2 \StoreAddress_reg[13]  ( .D(\add_60/A[13] ), .CK(clock), .RN(n412), 
        .Q(StoreAddress[13]) );
  DFFR_X2 \StoreAddress_reg[12]  ( .D(\add_60/A[12] ), .CK(clock), .RN(n412), 
        .Q(StoreAddress[12]) );
  DFFR_X2 \StoreAddress_reg[11]  ( .D(\add_60/A[11] ), .CK(clock), .RN(n412), 
        .Q(StoreAddress[11]) );
  DFFR_X2 \StoreAddress_reg[9]  ( .D(\add_60/A[9] ), .CK(clock), .RN(n411), 
        .Q(StoreAddress[9]) );
  DFFR_X2 \StoreAddress_reg[7]  ( .D(\add_60/A[7] ), .CK(clock), .RN(n411), 
        .Q(StoreAddress[7]) );
  DFFR_X2 \StoreAddress_reg[3]  ( .D(\add_60/A[3] ), .CK(clock), .RN(n410), 
        .Q(StoreAddress[3]) );
  DFFR_X2 \StoreAddress_reg[4]  ( .D(\add_60/A[4] ), .CK(clock), .RN(n410), 
        .Q(StoreAddress[4]) );
  DFFR_X2 \StoreAddress_reg[8]  ( .D(\add_60/A[8] ), .CK(clock), .RN(n411), 
        .Q(StoreAddress[8]) );
  DFFR_X2 \StoreAddress_reg[6]  ( .D(\add_60/A[6] ), .CK(clock), .RN(n411), 
        .Q(StoreAddress[6]) );
  DFFR_X2 \StoreAddress_reg[14]  ( .D(\add_60/A[14] ), .CK(clock), .RN(n412), 
        .Q(StoreAddress[14]) );
  DFFR_X2 \ReadAddress_reg[6]  ( .D(\U5/Z_6 ), .CK(clock), .RN(n411), .Q(
        \add_60/A[6] ) );
  DFFR_X2 \ReadAddress_reg[8]  ( .D(\U5/Z_8 ), .CK(clock), .RN(n411), .Q(
        \add_60/A[8] ) );
  DFFR_X2 \ReadAddress_reg[14]  ( .D(\U5/Z_14 ), .CK(clock), .RN(n412), .Q(
        \add_60/A[14] ), .QN(n442) );
  DFFR_X2 \AccumlateOut_reg[19]  ( .D(\U7/Z_19 ), .CK(clock), .RN(n413), .Q(
        AccumlateOut[19]) );
  DFFR_X2 \AccumlateOut_reg[18]  ( .D(\U7/Z_18 ), .CK(clock), .RN(n413), .Q(
        AccumlateOut[18]) );
  DFFR_X2 \AccumlateOut_reg[17]  ( .D(\U7/Z_17 ), .CK(clock), .RN(n413), .Q(
        AccumlateOut[17]) );
  DFFR_X2 \AccumlateOut_reg[16]  ( .D(\U7/Z_16 ), .CK(clock), .RN(n413), .Q(
        AccumlateOut[16]) );
  DFFR_X2 \AccumlateOut_reg[15]  ( .D(\U7/Z_15 ), .CK(clock), .RN(n413), .Q(
        AccumlateOut[15]) );
  DFFR_X2 \AccumlateOut_reg[14]  ( .D(\U7/Z_14 ), .CK(clock), .RN(n413), .Q(
        AccumlateOut[14]) );
  DFFR_X2 \AccumlateOut_reg[13]  ( .D(\U7/Z_13 ), .CK(clock), .RN(n414), .Q(
        AccumlateOut[13]) );
  DFFR_X2 \AccumlateOut_reg[12]  ( .D(\U7/Z_12 ), .CK(clock), .RN(n414), .Q(
        AccumlateOut[12]) );
  DFFR_X2 \AccumlateOut_reg[11]  ( .D(\U7/Z_11 ), .CK(clock), .RN(n414), .Q(
        AccumlateOut[11]) );
  DFFR_X2 \AccumlateOut_reg[10]  ( .D(\U7/Z_10 ), .CK(clock), .RN(n414), .Q(
        AccumlateOut[10]) );
  DFFR_X2 \AccumlateOut_reg[9]  ( .D(\U7/Z_9 ), .CK(clock), .RN(n414), .Q(
        AccumlateOut[9]) );
  DFFR_X2 \AccumlateOut_reg[4]  ( .D(\U7/Z_4 ), .CK(clock), .RN(n414), .Q(
        AccumlateOut[4]) );
  DFFR_X2 \AccumlateOut_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .RN(n414), .Q(
        AccumlateOut[3]) );
  NAND2_X2 U4 ( .A1(\add_60/A[4] ), .A2(n388), .ZN(n424) );
  AND4_X4 U6 ( .A1(n16), .A2(n17), .A3(n14), .A4(n15), .ZN(n375) );
  AND2_X1 U8 ( .A1(n1), .A2(start), .ZN(n376) );
  AND2_X1 U10 ( .A1(\add_63/A[8] ), .A2(start), .ZN(n377) );
  INV_X2 U12 ( .A(n379), .ZN(AccumlateOut[7]) );
  NOR2_X2 U14 ( .A1(n443), .A2(n442), .ZN(n444) );
  NAND2_X2 U16 ( .A1(n385), .A2(n392), .ZN(n422) );
  NAND2_X2 U17 ( .A1(\add_60/A[8] ), .A2(n389), .ZN(n432) );
  INV_X4 U20 ( .A(n381), .ZN(AccumlateOut[5]) );
  INV_X4 U21 ( .A(n383), .ZN(AccumlateOut[6]) );
  OR2_X4 U22 ( .A1(n402), .A2(n434), .ZN(n436) );
  INV_X2 U23 ( .A(n430), .ZN(n389) );
  OR2_X4 U24 ( .A1(n403), .A2(n436), .ZN(n438) );
  OR2_X4 U25 ( .A1(n390), .A2(n391), .ZN(n440) );
  OR2_X2 U26 ( .A1(n434), .A2(n402), .ZN(n390) );
  INV_X4 U27 ( .A(n422), .ZN(n388) );
  INV_X1 U28 ( .A(n385), .ZN(n418) );
  NOR2_X2 U29 ( .A1(n386), .A2(n33), .ZN(n385) );
  NOR2_X2 U36 ( .A1(n399), .A2(n424), .ZN(n387) );
  NAND2_X2 U37 ( .A1(\add_60/A[6] ), .A2(n387), .ZN(n428) );
  OR2_X1 U38 ( .A1(n404), .A2(n403), .ZN(n391) );
  NOR2_X2 U39 ( .A1(n397), .A2(n398), .ZN(n392) );
  NAND2_X2 U40 ( .A1(n34), .A2(n394), .ZN(n395) );
  NAND2_X1 U41 ( .A1(n393), .A2(n444), .ZN(n396) );
  NAND2_X2 U42 ( .A1(n395), .A2(n396), .ZN(n446) );
  INV_X2 U52 ( .A(n444), .ZN(n394) );
  INV_X4 U53 ( .A(n415), .ZN(n414) );
  INV_X4 U54 ( .A(n415), .ZN(n413) );
  INV_X4 U55 ( .A(n415), .ZN(n411) );
  INV_X4 U56 ( .A(n415), .ZN(n410) );
  INV_X4 U57 ( .A(n415), .ZN(n412) );
  INV_X4 U58 ( .A(reset_n), .ZN(n415) );
  OAI21_X2 U59 ( .B1(n11), .B2(n2), .A(n4), .ZN(n48) );
  OR2_X1 U60 ( .A1(n397), .A2(n418), .ZN(n420) );
  OR2_X1 U61 ( .A1(n399), .A2(n424), .ZN(n426) );
  OR2_X1 U62 ( .A1(n400), .A2(n428), .ZN(n430) );
  OR2_X1 U63 ( .A1(n401), .A2(n432), .ZN(n434) );
  OR2_X1 U64 ( .A1(n405), .A2(n440), .ZN(n443) );
  INV_X2 U65 ( .A(n406), .ZN(AccumlateOut[0]) );
  INV_X2 U66 ( .A(n408), .ZN(AccumlateOut[1]) );
  INV_X4 U67 ( .A(start), .ZN(n36) );
  NAND2_X2 U68 ( .A1(n2), .A2(start), .ZN(n4) );
  NAND2_X2 U69 ( .A1(start), .A2(n1), .ZN(n2) );
  NOR2_X2 U70 ( .A1(\add_60/A[0] ), .A2(n2), .ZN(\U5/Z_0 ) );
  XNOR2_X2 U71 ( .A(\add_60/A[0] ), .B(\add_60/A[1] ), .ZN(n416) );
  NOR2_X2 U72 ( .A1(n2), .A2(n416), .ZN(\U5/Z_1 ) );
  XOR2_X2 U73 ( .A(n418), .B(\add_60/A[2] ), .Z(n417) );
  NOR2_X2 U74 ( .A1(n2), .A2(n417), .ZN(\U5/Z_2 ) );
  XOR2_X2 U75 ( .A(n420), .B(\add_60/A[3] ), .Z(n419) );
  NOR2_X2 U76 ( .A1(n2), .A2(n419), .ZN(\U5/Z_3 ) );
  XOR2_X2 U77 ( .A(n422), .B(\add_60/A[4] ), .Z(n421) );
  NOR2_X2 U78 ( .A1(n2), .A2(n421), .ZN(\U5/Z_4 ) );
  XOR2_X2 U79 ( .A(n424), .B(\add_60/A[5] ), .Z(n423) );
  NOR2_X2 U80 ( .A1(n2), .A2(n423), .ZN(\U5/Z_5 ) );
  XOR2_X2 U81 ( .A(n426), .B(\add_60/A[6] ), .Z(n425) );
  NOR2_X2 U82 ( .A1(n2), .A2(n425), .ZN(\U5/Z_6 ) );
  XOR2_X2 U83 ( .A(n428), .B(\add_60/A[7] ), .Z(n427) );
  NOR2_X2 U84 ( .A1(n2), .A2(n427), .ZN(\U5/Z_7 ) );
  XOR2_X2 U85 ( .A(n430), .B(\add_60/A[8] ), .Z(n429) );
  NOR2_X2 U86 ( .A1(n2), .A2(n429), .ZN(\U5/Z_8 ) );
  XOR2_X2 U87 ( .A(n432), .B(\add_60/A[9] ), .Z(n431) );
  NOR2_X2 U88 ( .A1(n2), .A2(n431), .ZN(\U5/Z_9 ) );
  XOR2_X2 U89 ( .A(n434), .B(\add_60/A[10] ), .Z(n433) );
  NOR2_X2 U90 ( .A1(n2), .A2(n433), .ZN(\U5/Z_10 ) );
  XOR2_X2 U91 ( .A(n436), .B(\add_60/A[11] ), .Z(n435) );
  NOR2_X2 U92 ( .A1(n2), .A2(n435), .ZN(\U5/Z_11 ) );
  XOR2_X2 U93 ( .A(n438), .B(\add_60/A[12] ), .Z(n437) );
  NOR2_X2 U94 ( .A1(n2), .A2(n437), .ZN(\U5/Z_12 ) );
  XOR2_X2 U95 ( .A(n440), .B(\add_60/A[13] ), .Z(n439) );
  NOR2_X2 U96 ( .A1(n2), .A2(n439), .ZN(\U5/Z_13 ) );
  XOR2_X2 U97 ( .A(n443), .B(\add_60/A[14] ), .Z(n441) );
  NOR2_X2 U98 ( .A1(n2), .A2(n441), .ZN(\U5/Z_14 ) );
  INV_X4 U99 ( .A(\U4/DATA3_0 ), .ZN(n445) );
  OAI22_X2 U100 ( .A1(n2), .A2(n446), .B1(start), .B2(n445), .ZN(\U4/Z_0 ) );
  AND2_X1 U101 ( .A1(\U8/DATA1_0 ), .A2(n375), .ZN(\U7/Z_0 ) );
  AND2_X1 U102 ( .A1(\U8/DATA1_1 ), .A2(n375), .ZN(\U7/Z_1 ) );
  AND2_X1 U103 ( .A1(\U8/DATA1_2 ), .A2(n375), .ZN(\U7/Z_2 ) );
  AND2_X1 U104 ( .A1(\U8/DATA1_3 ), .A2(n375), .ZN(\U7/Z_3 ) );
  AND2_X1 U105 ( .A1(\U8/DATA1_4 ), .A2(n375), .ZN(\U7/Z_4 ) );
  AND2_X1 U106 ( .A1(\U8/DATA1_5 ), .A2(n375), .ZN(\U7/Z_5 ) );
  AND2_X1 U107 ( .A1(\U8/DATA1_6 ), .A2(n375), .ZN(\U7/Z_6 ) );
  AND2_X1 U108 ( .A1(\U8/DATA1_7 ), .A2(n375), .ZN(\U7/Z_7 ) );
  AND2_X1 U109 ( .A1(\U8/DATA1_8 ), .A2(n375), .ZN(\U7/Z_8 ) );
  AND2_X1 U110 ( .A1(\U8/DATA1_9 ), .A2(n375), .ZN(\U7/Z_9 ) );
  AND2_X1 U111 ( .A1(\U8/DATA1_10 ), .A2(n375), .ZN(\U7/Z_10 ) );
  AND2_X1 U112 ( .A1(\U8/DATA1_11 ), .A2(n375), .ZN(\U7/Z_11 ) );
  AND2_X1 U113 ( .A1(\U8/DATA1_12 ), .A2(n375), .ZN(\U7/Z_12 ) );
  AND2_X1 U114 ( .A1(\U8/DATA1_13 ), .A2(n375), .ZN(\U7/Z_13 ) );
  INV_X4 U115 ( .A(\U3/U1/DATA1_7 ), .ZN(n10) );
  INV_X4 U116 ( .A(\U3/U1/DATA1_6 ), .ZN(n9) );
  INV_X4 U117 ( .A(\U3/U1/DATA1_5 ), .ZN(n8) );
  INV_X4 U118 ( .A(\U3/U1/DATA1_4 ), .ZN(n7) );
  INV_X4 U119 ( .A(\U3/U1/DATA1_3 ), .ZN(n6) );
  INV_X4 U120 ( .A(\U3/U1/DATA1_2 ), .ZN(n5) );
  INV_X4 U121 ( .A(\U3/U1/DATA1_1 ), .ZN(n3) );
endmodule


module Cdf_Accumlate ( clock, reset_n, AccumlateIn, StartIn, StoreAddressIn, 
        AccumlateResult, StoreAddressOut, StartOut, CdfMin, CdfValid );
  input [19:0] AccumlateIn;
  input [15:0] StoreAddressIn;
  output [19:0] AccumlateResult;
  output [15:0] StoreAddressOut;
  output [19:0] CdfMin;
  input clock, reset_n, StartIn;
  output StartOut, CdfValid;
  wire   \U8/Z_0 , \U6/DATA2_0 , \U6/DATA2_1 , \U6/DATA2_2 , \U6/DATA2_3 ,
         \U6/DATA2_4 , \U6/DATA2_5 , \U6/DATA2_6 , \U6/DATA2_7 , \U6/DATA2_8 ,
         \U6/DATA2_9 , \U6/DATA2_10 , \U6/DATA2_11 , \U6/DATA2_12 ,
         \U6/DATA2_13 , \U6/DATA2_14 , \U6/DATA2_15 , \U6/DATA2_16 ,
         \U6/DATA2_17 , \U6/DATA2_18 , \U6/DATA2_19 , \add/B[0] , \add/B[1] ,
         \add/B[2] , \add/B[3] , \add/B[4] , \add/B[5] , \add/B[6] ,
         \add/B[7] , \add/B[8] , \add/B[9] , \add/B[10] , \add/B[11] ,
         \add/B[12] , \add/B[13] , \add/B[14] , \add/B[15] , \add/B[16] ,
         \add/B[17] , \add/B[18] , \add/B[19] , \add/A[0] , \add/A[1] ,
         \add/A[2] , \add/A[3] , \add/A[4] , \add/A[5] , \add/A[6] ,
         \add/A[7] , \add/A[8] , \add/A[9] , \add/A[10] , \add/A[11] ,
         \add/A[12] , \add/A[13] , \add/A[14] , \add/A[15] , \add/A[16] ,
         \add/A[17] , \add/A[18] , \add/A[19] , n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n64, n65, n79, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459;
  assign CdfMin[0] = \U6/DATA2_0 ;
  assign CdfMin[1] = \U6/DATA2_1 ;
  assign CdfMin[2] = \U6/DATA2_2 ;
  assign CdfMin[3] = \U6/DATA2_3 ;
  assign CdfMin[4] = \U6/DATA2_4 ;
  assign CdfMin[5] = \U6/DATA2_5 ;
  assign CdfMin[6] = \U6/DATA2_6 ;
  assign CdfMin[7] = \U6/DATA2_7 ;
  assign CdfMin[8] = \U6/DATA2_8 ;
  assign CdfMin[9] = \U6/DATA2_9 ;
  assign CdfMin[10] = \U6/DATA2_10 ;
  assign CdfMin[11] = \U6/DATA2_11 ;
  assign CdfMin[12] = \U6/DATA2_12 ;
  assign CdfMin[13] = \U6/DATA2_13 ;
  assign CdfMin[14] = \U6/DATA2_14 ;
  assign CdfMin[15] = \U6/DATA2_15 ;
  assign CdfMin[16] = \U6/DATA2_16 ;
  assign CdfMin[17] = \U6/DATA2_17 ;
  assign CdfMin[18] = \U6/DATA2_18 ;
  assign CdfMin[19] = \U6/DATA2_19 ;
  assign \add/B[0]  = AccumlateIn[0];
  assign \add/B[1]  = AccumlateIn[1];
  assign \add/B[2]  = AccumlateIn[2];
  assign \add/B[3]  = AccumlateIn[3];
  assign \add/B[4]  = AccumlateIn[4];
  assign \add/B[5]  = AccumlateIn[5];
  assign \add/B[6]  = AccumlateIn[6];
  assign \add/B[7]  = AccumlateIn[7];
  assign \add/B[8]  = AccumlateIn[8];
  assign \add/B[9]  = AccumlateIn[9];
  assign \add/B[10]  = AccumlateIn[10];
  assign \add/B[11]  = AccumlateIn[11];
  assign \add/B[12]  = AccumlateIn[12];
  assign \add/B[13]  = AccumlateIn[13];
  assign \add/B[14]  = AccumlateIn[14];
  assign \add/B[15]  = AccumlateIn[15];
  assign \add/B[16]  = AccumlateIn[16];
  assign \add/B[17]  = AccumlateIn[17];
  assign \add/B[18]  = AccumlateIn[18];
  assign \add/B[19]  = AccumlateIn[19];
  assign AccumlateResult[0] = \add/A[0] ;
  assign AccumlateResult[1] = \add/A[1] ;
  assign AccumlateResult[2] = \add/A[2] ;
  assign AccumlateResult[3] = \add/A[3] ;
  assign AccumlateResult[4] = \add/A[4] ;
  assign AccumlateResult[5] = \add/A[5] ;
  assign AccumlateResult[6] = \add/A[6] ;
  assign AccumlateResult[7] = \add/A[7] ;
  assign AccumlateResult[8] = \add/A[8] ;
  assign AccumlateResult[9] = \add/A[9] ;
  assign AccumlateResult[10] = \add/A[10] ;
  assign AccumlateResult[11] = \add/A[11] ;
  assign AccumlateResult[12] = \add/A[12] ;
  assign AccumlateResult[13] = \add/A[13] ;
  assign AccumlateResult[14] = \add/A[14] ;
  assign AccumlateResult[15] = \add/A[15] ;
  assign AccumlateResult[16] = \add/A[16] ;
  assign AccumlateResult[17] = \add/A[17] ;
  assign AccumlateResult[18] = \add/A[18] ;
  assign AccumlateResult[19] = \add/A[19] ;

  DFF_X1 \StoreAddressOut_reg[15]  ( .D(StoreAddressIn[15]), .CK(clock), .Q(
        StoreAddressOut[15]) );
  DFF_X1 \StoreAddressOut_reg[14]  ( .D(StoreAddressIn[14]), .CK(clock), .Q(
        StoreAddressOut[14]) );
  DFF_X1 \StoreAddressOut_reg[13]  ( .D(StoreAddressIn[13]), .CK(clock), .Q(
        StoreAddressOut[13]) );
  DFF_X1 \StoreAddressOut_reg[12]  ( .D(StoreAddressIn[12]), .CK(clock), .Q(
        StoreAddressOut[12]) );
  DFF_X1 \StoreAddressOut_reg[11]  ( .D(StoreAddressIn[11]), .CK(clock), .Q(
        StoreAddressOut[11]) );
  DFF_X1 \StoreAddressOut_reg[10]  ( .D(StoreAddressIn[10]), .CK(clock), .Q(
        StoreAddressOut[10]) );
  DFF_X1 \StoreAddressOut_reg[9]  ( .D(StoreAddressIn[9]), .CK(clock), .Q(
        StoreAddressOut[9]) );
  DFF_X1 \StoreAddressOut_reg[8]  ( .D(StoreAddressIn[8]), .CK(clock), .Q(
        StoreAddressOut[8]) );
  DFF_X1 \StoreAddressOut_reg[7]  ( .D(StoreAddressIn[7]), .CK(clock), .Q(
        StoreAddressOut[7]) );
  DFF_X1 \StoreAddressOut_reg[6]  ( .D(StoreAddressIn[6]), .CK(clock), .Q(
        StoreAddressOut[6]) );
  DFF_X1 \StoreAddressOut_reg[5]  ( .D(StoreAddressIn[5]), .CK(clock), .Q(
        StoreAddressOut[5]) );
  DFF_X1 \StoreAddressOut_reg[4]  ( .D(StoreAddressIn[4]), .CK(clock), .Q(
        StoreAddressOut[4]) );
  DFF_X1 \StoreAddressOut_reg[3]  ( .D(StoreAddressIn[3]), .CK(clock), .Q(
        StoreAddressOut[3]) );
  DFF_X1 \StoreAddressOut_reg[2]  ( .D(StoreAddressIn[2]), .CK(clock), .Q(
        StoreAddressOut[2]) );
  DFF_X1 \StoreAddressOut_reg[1]  ( .D(StoreAddressIn[1]), .CK(clock), .Q(
        StoreAddressOut[1]) );
  DFF_X1 \StoreAddressOut_reg[0]  ( .D(StoreAddressIn[0]), .CK(clock), .Q(
        StoreAddressOut[0]) );
  AND3_X2 U25 ( .A1(n22), .A2(n64), .A3(StartIn), .ZN(\U8/Z_0 ) );
  NAND3_X2 U35 ( .A1(n38), .A2(n37), .A3(n39), .ZN(n79) );
  INV_X4 U80 ( .A(n65), .ZN(n22) );
  DFFR_X2 \AccumlateResult_reg[0]  ( .D(n459), .CK(clock), .RN(n264), .Q(
        \add/A[0] ), .QN(n253) );
  DFFR_X2 \AccumlateResult_reg[1]  ( .D(n458), .CK(clock), .RN(n264), .Q(
        \add/A[1] ), .QN(n252) );
  DFFR_X2 \AccumlateResult_reg[2]  ( .D(n457), .CK(clock), .RN(n264), .Q(
        \add/A[2] ), .QN(n245) );
  DFFR_X2 \AccumlateResult_reg[8]  ( .D(n451), .CK(clock), .RN(n263), .Q(
        \add/A[8] ), .QN(n242) );
  DFFR_X2 \AccumlateResult_reg[5]  ( .D(n454), .CK(clock), .RN(n263), .Q(
        \add/A[5] ), .QN(n241) );
  DFFR_X2 \AccumlateResult_reg[4]  ( .D(n455), .CK(clock), .RN(reset_n), .Q(
        \add/A[4] ), .QN(n318) );
  DFFR_X2 \CdfMin_reg[15]  ( .D(n86), .CK(clock), .RN(n264), .Q(\U6/DATA2_15 ), 
        .QN(n26) );
  DFFR_X2 \CdfMin_reg[17]  ( .D(n84), .CK(clock), .RN(n264), .Q(\U6/DATA2_17 ), 
        .QN(n24) );
  DFFR_X2 \CdfMin_reg[18]  ( .D(n83), .CK(clock), .RN(n264), .Q(\U6/DATA2_18 ), 
        .QN(n23) );
  DFFR_X2 \CdfMin_reg[14]  ( .D(n87), .CK(clock), .RN(n264), .Q(\U6/DATA2_14 ), 
        .QN(n27) );
  DFFR_X2 \CdfMin_reg[3]  ( .D(n98), .CK(clock), .RN(n262), .Q(\U6/DATA2_3 ), 
        .QN(n38) );
  DFFR_X2 \CdfMin_reg[8]  ( .D(n93), .CK(clock), .RN(n262), .Q(\U6/DATA2_8 ), 
        .QN(n33) );
  DFFR_X2 \CdfMin_reg[7]  ( .D(n94), .CK(clock), .RN(n262), .Q(\U6/DATA2_7 ), 
        .QN(n34) );
  DFFR_X2 \CdfMin_reg[10]  ( .D(n91), .CK(clock), .RN(n262), .Q(\U6/DATA2_10 ), 
        .QN(n31) );
  DFFR_X2 \CdfMin_reg[9]  ( .D(n92), .CK(clock), .RN(n262), .Q(\U6/DATA2_9 ), 
        .QN(n32) );
  DFFR_X2 \CdfMin_reg[12]  ( .D(n89), .CK(clock), .RN(n262), .Q(\U6/DATA2_12 ), 
        .QN(n29) );
  DFFR_X2 \CdfMin_reg[11]  ( .D(n90), .CK(clock), .RN(n262), .Q(\U6/DATA2_11 ), 
        .QN(n30) );
  DFFR_X2 \CdfMin_reg[2]  ( .D(n99), .CK(clock), .RN(n262), .Q(\U6/DATA2_2 ), 
        .QN(n39) );
  DFFR_X2 \CdfMin_reg[4]  ( .D(n97), .CK(clock), .RN(n262), .Q(\U6/DATA2_4 ), 
        .QN(n37) );
  DFFR_X2 \CdfMin_reg[1]  ( .D(n100), .CK(clock), .RN(n262), .Q(\U6/DATA2_1 ), 
        .QN(n40) );
  DFFR_X2 \CdfMin_reg[5]  ( .D(n96), .CK(clock), .RN(n262), .Q(\U6/DATA2_5 ), 
        .QN(n36) );
  DFFR_X2 \CdfMin_reg[0]  ( .D(n101), .CK(clock), .RN(n264), .Q(\U6/DATA2_0 ), 
        .QN(n41) );
  DFFR_X2 \CdfMin_reg[13]  ( .D(n88), .CK(clock), .RN(n264), .Q(\U6/DATA2_13 ), 
        .QN(n28) );
  DFFR_X2 \CdfMin_reg[6]  ( .D(n95), .CK(clock), .RN(n262), .Q(\U6/DATA2_6 ), 
        .QN(n35) );
  DFFR_X2 \CdfMin_reg[19]  ( .D(n82), .CK(clock), .RN(reset_n), .Q(
        \U6/DATA2_19 ), .QN(n21) );
  DFFR_X2 \CdfMin_reg[16]  ( .D(n85), .CK(clock), .RN(n264), .Q(\U6/DATA2_16 ), 
        .QN(n25) );
  DFFR_X2 \AccumlateResult_reg[6]  ( .D(n453), .CK(clock), .RN(n263), .Q(
        \add/A[6] ), .QN(n230) );
  DFFR_X2 \AccumlateResult_reg[7]  ( .D(n452), .CK(clock), .RN(n263), .Q(
        \add/A[7] ), .QN(n251) );
  DFFR_X2 \AccumlateResult_reg[10]  ( .D(n449), .CK(clock), .RN(n263), .Q(
        \add/A[10] ), .QN(n379) );
  DFFR_X2 \AccumlateResult_reg[13]  ( .D(n446), .CK(clock), .RN(n263), .Q(
        \add/A[13] ), .QN(n385) );
  DFFR_X2 \AccumlateResult_reg[3]  ( .D(n456), .CK(clock), .RN(n264), .Q(
        \add/A[3] ), .QN(n381) );
  DFFR_X2 CdfValid_reg ( .D(\U8/Z_0 ), .CK(clock), .RN(reset_n), .Q(CdfValid)
         );
  DFFR_X2 \AccumlateResult_reg[16]  ( .D(n443), .CK(clock), .RN(n263), .Q(
        \add/A[16] ) );
  DFFR_X2 StartOut_reg ( .D(StartIn), .CK(clock), .RN(n264), .Q(StartOut) );
  DFFR_X2 \AccumlateResult_reg[9]  ( .D(n450), .CK(clock), .RN(n263), .Q(
        \add/A[9] ), .QN(n380) );
  DFFR_X2 \AccumlateResult_reg[12]  ( .D(n447), .CK(clock), .RN(n263), .Q(
        \add/A[12] ), .QN(n273) );
  DFFR_X2 \AccumlateResult_reg[11]  ( .D(n448), .CK(clock), .RN(n263), .Q(
        \add/A[11] ), .QN(n386) );
  DFFR_X2 \AccumlateResult_reg[17]  ( .D(n442), .CK(clock), .RN(reset_n), .Q(
        \add/A[17] ), .QN(n406) );
  DFFR_X2 \AccumlateResult_reg[18]  ( .D(n441), .CK(clock), .RN(reset_n), .Q(
        \add/A[18] ), .QN(n423) );
  DFFR_X2 \AccumlateResult_reg[19]  ( .D(n440), .CK(clock), .RN(reset_n), .Q(
        \add/A[19] ), .QN(n419) );
  DFFR_X2 \AccumlateResult_reg[14]  ( .D(n445), .CK(clock), .RN(n263), .Q(
        \add/A[14] ), .QN(n270) );
  DFFR_X2 \AccumlateResult_reg[15]  ( .D(n444), .CK(clock), .RN(n263), .Q(
        \add/A[15] ), .QN(n268) );
  AND2_X2 U3 ( .A1(n330), .A2(n335), .ZN(n216) );
  AOI22_X4 U4 ( .A1(n297), .A2(n224), .B1(\add/B[11] ), .B2(\add/A[11] ), .ZN(
        n359) );
  INV_X1 U5 ( .A(n287), .ZN(n275) );
  INV_X2 U6 ( .A(n292), .ZN(n288) );
  OAI21_X2 U7 ( .B1(n369), .B2(n304), .A(n303), .ZN(n425) );
  AOI22_X4 U8 ( .A1(n302), .A2(n301), .B1(\add/B[15] ), .B2(\add/A[15] ), .ZN(
        n369) );
  AOI22_X4 U9 ( .A1(n298), .A2(n299), .B1(\add/B[12] ), .B2(\add/A[12] ), .ZN(
        n362) );
  NAND3_X2 U10 ( .A1(n327), .A2(n329), .A3(n288), .ZN(n293) );
  NAND2_X2 U11 ( .A1(n241), .A2(n289), .ZN(n329) );
  AOI221_X2 U12 ( .B1(n238), .B2(n379), .C1(n240), .C2(n347), .A(n239), .ZN(
        n237) );
  OAI22_X2 U13 ( .A1(n362), .A2(n229), .B1(n271), .B2(n385), .ZN(n228) );
  NAND2_X2 U14 ( .A1(n246), .A2(n287), .ZN(n292) );
  XNOR2_X1 U15 ( .A(n360), .B(n298), .ZN(n361) );
  AND2_X2 U16 ( .A1(\add/B[0] ), .A2(n254), .ZN(n219) );
  AND2_X1 U17 ( .A1(n296), .A2(n295), .ZN(n221) );
  NAND3_X1 U18 ( .A1(n253), .A2(n419), .A3(n384), .ZN(n388) );
  OAI22_X2 U19 ( .A1(n226), .A2(n229), .B1(n271), .B2(n385), .ZN(n227) );
  INV_X2 U20 ( .A(n225), .ZN(n226) );
  NOR3_X1 U21 ( .A1(n217), .A2(n222), .A3(n429), .ZN(n430) );
  INV_X1 U22 ( .A(n392), .ZN(n443) );
  AOI22_X4 U23 ( .A1(n228), .A2(n300), .B1(\add/B[14] ), .B2(\add/A[14] ), 
        .ZN(n366) );
  AND2_X2 U24 ( .A1(n428), .A2(n427), .ZN(n217) );
  AND2_X4 U26 ( .A1(n429), .A2(n424), .ZN(n218) );
  AND2_X4 U27 ( .A1(n307), .A2(n308), .ZN(n220) );
  AND2_X4 U28 ( .A1(n423), .A2(n422), .ZN(n222) );
  AND2_X4 U29 ( .A1(StartIn), .A2(n432), .ZN(n223) );
  XOR2_X1 U30 ( .A(n318), .B(\add/B[4] ), .Z(n320) );
  INV_X2 U31 ( .A(\add/B[4] ), .ZN(n285) );
  INV_X4 U32 ( .A(n369), .ZN(n370) );
  NAND2_X2 U33 ( .A1(n223), .A2(n431), .ZN(n433) );
  NOR3_X2 U34 ( .A1(n232), .A2(n233), .A3(n430), .ZN(n431) );
  NAND2_X2 U36 ( .A1(n296), .A2(n295), .ZN(n224) );
  NAND2_X2 U37 ( .A1(n220), .A2(n313), .ZN(n281) );
  INV_X1 U38 ( .A(n362), .ZN(n225) );
  AND2_X4 U39 ( .A1(n385), .A2(n271), .ZN(n229) );
  NOR4_X1 U40 ( .A1(\U6/DATA2_0 ), .A2(\U6/DATA2_19 ), .A3(\U6/DATA2_18 ), 
        .A4(\U6/DATA2_14 ), .ZN(n376) );
  XNOR2_X1 U41 ( .A(\add/B[8] ), .B(\add/A[8] ), .ZN(n236) );
  XNOR2_X1 U42 ( .A(n219), .B(n231), .ZN(n306) );
  XOR2_X1 U43 ( .A(n278), .B(\add/A[1] ), .Z(n231) );
  XOR2_X1 U44 ( .A(\add/B[0] ), .B(\add/A[0] ), .Z(n266) );
  AND2_X1 U45 ( .A1(n222), .A2(n218), .ZN(n232) );
  AND2_X2 U46 ( .A1(n217), .A2(n218), .ZN(n233) );
  INV_X4 U47 ( .A(n265), .ZN(n263) );
  INV_X4 U48 ( .A(n265), .ZN(n264) );
  INV_X4 U49 ( .A(n265), .ZN(n262) );
  INV_X4 U50 ( .A(reset_n), .ZN(n265) );
  INV_X4 U51 ( .A(n248), .ZN(n308) );
  INV_X4 U52 ( .A(n350), .ZN(n239) );
  NAND2_X2 U53 ( .A1(n257), .A2(n64), .ZN(n439) );
  NAND2_X2 U54 ( .A1(n437), .A2(n64), .ZN(n259) );
  OR2_X1 U55 ( .A1(n244), .A2(n234), .ZN(n342) );
  AND2_X4 U56 ( .A1(n216), .A2(n340), .ZN(n234) );
  OR2_X1 U57 ( .A1(\add/A[11] ), .A2(\add/B[11] ), .ZN(n297) );
  XNOR2_X2 U58 ( .A(n235), .B(n407), .ZN(n305) );
  XNOR2_X2 U59 ( .A(n406), .B(\add/B[17] ), .ZN(n235) );
  INV_X4 U60 ( .A(\add/B[10] ), .ZN(n238) );
  XNOR2_X2 U61 ( .A(n343), .B(n236), .ZN(n344) );
  INV_X4 U62 ( .A(StartIn), .ZN(n260) );
  NAND2_X1 U63 ( .A1(n347), .A2(n346), .ZN(n351) );
  INV_X4 U64 ( .A(n237), .ZN(n295) );
  AND2_X4 U65 ( .A1(n346), .A2(n352), .ZN(n240) );
  INV_X4 U66 ( .A(n345), .ZN(n347) );
  INV_X4 U67 ( .A(n333), .ZN(n243) );
  NAND2_X1 U68 ( .A1(\add/B[3] ), .A2(\add/A[3] ), .ZN(n284) );
  XOR2_X1 U69 ( .A(\add/B[3] ), .B(\add/A[3] ), .Z(n315) );
  XNOR2_X1 U70 ( .A(\add/B[2] ), .B(\add/A[2] ), .ZN(n309) );
  INV_X1 U71 ( .A(n246), .ZN(n244) );
  NAND2_X1 U72 ( .A1(n312), .A2(n311), .ZN(n314) );
  NAND2_X1 U73 ( .A1(n330), .A2(n340), .ZN(n334) );
  INV_X4 U74 ( .A(\add/B[1] ), .ZN(n278) );
  NOR2_X2 U75 ( .A1(n243), .A2(n247), .ZN(n246) );
  AND2_X4 U76 ( .A1(n251), .A2(n250), .ZN(n247) );
  INV_X2 U77 ( .A(n255), .ZN(n256) );
  NOR2_X2 U78 ( .A1(n278), .A2(n252), .ZN(n248) );
  NOR4_X1 U79 ( .A1(n383), .A2(n382), .A3(\add/A[4] ), .A4(\add/A[5] ), .ZN(
        n390) );
  XOR2_X1 U81 ( .A(\add/B[5] ), .B(\add/A[5] ), .Z(n324) );
  NAND2_X1 U82 ( .A1(n219), .A2(n279), .ZN(n249) );
  INV_X1 U83 ( .A(\add/B[7] ), .ZN(n250) );
  NAND2_X1 U84 ( .A1(\add/B[6] ), .A2(\add/A[6] ), .ZN(n335) );
  XOR2_X1 U85 ( .A(\add/B[6] ), .B(\add/A[6] ), .Z(n331) );
  NAND2_X2 U86 ( .A1(n219), .A2(n279), .ZN(n307) );
  INV_X2 U87 ( .A(n253), .ZN(n254) );
  NAND2_X2 U88 ( .A1(n282), .A2(n311), .ZN(n255) );
  NAND2_X2 U89 ( .A1(n256), .A2(n281), .ZN(n283) );
  NAND2_X1 U90 ( .A1(n308), .A2(n249), .ZN(n312) );
  NAND2_X1 U91 ( .A1(n327), .A2(n328), .ZN(n323) );
  NOR3_X1 U92 ( .A1(\add/A[8] ), .A2(\add/A[7] ), .A3(\add/A[6] ), .ZN(n378)
         );
  XOR2_X1 U93 ( .A(\add/B[7] ), .B(\add/A[7] ), .Z(n337) );
  NAND2_X1 U94 ( .A1(\add/B[7] ), .A2(\add/A[7] ), .ZN(n341) );
  INV_X1 U95 ( .A(n433), .ZN(n440) );
  NAND3_X1 U96 ( .A1(n329), .A2(n328), .A3(n327), .ZN(n340) );
  INV_X1 U97 ( .A(n366), .ZN(n367) );
  INV_X1 U98 ( .A(n425), .ZN(n407) );
  NOR3_X1 U99 ( .A1(n410), .A2(n409), .A3(n425), .ZN(n411) );
  NAND2_X2 U100 ( .A1(StartIn), .A2(n65), .ZN(n257) );
  NAND2_X2 U101 ( .A1(StartIn), .A2(n65), .ZN(n258) );
  NAND2_X2 U102 ( .A1(StartIn), .A2(n266), .ZN(n434) );
  INV_X4 U103 ( .A(n434), .ZN(n459) );
  INV_X4 U104 ( .A(\add/B[15] ), .ZN(n267) );
  NAND2_X2 U105 ( .A1(n268), .A2(n267), .ZN(n302) );
  INV_X4 U106 ( .A(\add/B[14] ), .ZN(n269) );
  NAND2_X2 U107 ( .A1(n270), .A2(n269), .ZN(n300) );
  INV_X4 U108 ( .A(\add/B[13] ), .ZN(n271) );
  INV_X4 U109 ( .A(\add/B[12] ), .ZN(n272) );
  NAND2_X2 U110 ( .A1(n273), .A2(n272), .ZN(n299) );
  NAND2_X2 U111 ( .A1(\add/B[10] ), .A2(\add/A[10] ), .ZN(n296) );
  INV_X4 U112 ( .A(\add/B[8] ), .ZN(n274) );
  NAND2_X2 U113 ( .A1(n242), .A2(n274), .ZN(n287) );
  OAI22_X2 U114 ( .A1(n275), .A2(n341), .B1(n242), .B2(n274), .ZN(n276) );
  INV_X4 U115 ( .A(n276), .ZN(n346) );
  NAND2_X2 U116 ( .A1(\add/B[9] ), .A2(\add/A[9] ), .ZN(n352) );
  INV_X4 U117 ( .A(\add/B[3] ), .ZN(n277) );
  NAND2_X2 U118 ( .A1(n381), .A2(n277), .ZN(n282) );
  NAND2_X2 U119 ( .A1(\add/B[2] ), .A2(\add/A[2] ), .ZN(n313) );
  NAND2_X2 U120 ( .A1(n252), .A2(n278), .ZN(n279) );
  INV_X4 U121 ( .A(\add/B[2] ), .ZN(n280) );
  NAND2_X2 U122 ( .A1(n245), .A2(n280), .ZN(n311) );
  NAND2_X2 U123 ( .A1(n283), .A2(n284), .ZN(n328) );
  INV_X4 U124 ( .A(n328), .ZN(n319) );
  NAND2_X2 U125 ( .A1(n318), .A2(n285), .ZN(n327) );
  INV_X4 U126 ( .A(\add/B[5] ), .ZN(n289) );
  INV_X4 U127 ( .A(\add/B[6] ), .ZN(n286) );
  NAND2_X2 U128 ( .A1(n230), .A2(n286), .ZN(n333) );
  INV_X4 U129 ( .A(n329), .ZN(n290) );
  NAND2_X2 U130 ( .A1(\add/B[4] ), .A2(\add/A[4] ), .ZN(n322) );
  OAI22_X2 U131 ( .A1(n290), .A2(n322), .B1(n241), .B2(n289), .ZN(n291) );
  INV_X4 U132 ( .A(n291), .ZN(n330) );
  OAI22_X2 U133 ( .A1(n319), .A2(n293), .B1(n216), .B2(n292), .ZN(n345) );
  INV_X4 U134 ( .A(\add/B[9] ), .ZN(n294) );
  NAND2_X2 U135 ( .A1(n380), .A2(n294), .ZN(n350) );
  INV_X4 U136 ( .A(n359), .ZN(n298) );
  INV_X4 U137 ( .A(n366), .ZN(n301) );
  NOR2_X2 U138 ( .A1(\add/B[16] ), .A2(\add/A[16] ), .ZN(n304) );
  NAND2_X2 U139 ( .A1(\add/B[16] ), .A2(\add/A[16] ), .ZN(n303) );
  NAND2_X2 U140 ( .A1(StartIn), .A2(n305), .ZN(n391) );
  INV_X4 U141 ( .A(n391), .ZN(n442) );
  NAND2_X2 U142 ( .A1(StartIn), .A2(n306), .ZN(n400) );
  INV_X4 U143 ( .A(n400), .ZN(n458) );
  XNOR2_X2 U144 ( .A(n309), .B(n312), .ZN(n310) );
  NAND2_X2 U145 ( .A1(StartIn), .A2(n310), .ZN(n435) );
  INV_X4 U146 ( .A(n435), .ZN(n457) );
  NAND2_X2 U147 ( .A1(n314), .A2(n313), .ZN(n316) );
  XOR2_X2 U148 ( .A(n316), .B(n315), .Z(n317) );
  NAND2_X2 U149 ( .A1(StartIn), .A2(n317), .ZN(n436) );
  INV_X4 U150 ( .A(n436), .ZN(n456) );
  XOR2_X2 U151 ( .A(n320), .B(n319), .Z(n321) );
  NAND2_X2 U152 ( .A1(StartIn), .A2(n321), .ZN(n438) );
  INV_X4 U153 ( .A(n438), .ZN(n455) );
  NAND2_X2 U154 ( .A1(n323), .A2(n322), .ZN(n325) );
  XOR2_X2 U155 ( .A(n325), .B(n324), .Z(n326) );
  NAND2_X2 U156 ( .A1(StartIn), .A2(n326), .ZN(n401) );
  INV_X4 U157 ( .A(n401), .ZN(n454) );
  XOR2_X2 U158 ( .A(n334), .B(n331), .Z(n332) );
  NAND2_X2 U159 ( .A1(StartIn), .A2(n332), .ZN(n402) );
  INV_X4 U160 ( .A(n402), .ZN(n453) );
  NAND2_X2 U161 ( .A1(n334), .A2(n333), .ZN(n336) );
  NAND2_X2 U162 ( .A1(n336), .A2(n335), .ZN(n338) );
  XOR2_X2 U163 ( .A(n338), .B(n337), .Z(n339) );
  NAND2_X2 U164 ( .A1(StartIn), .A2(n339), .ZN(n399) );
  INV_X4 U165 ( .A(n399), .ZN(n452) );
  NAND2_X2 U166 ( .A1(n342), .A2(n341), .ZN(n343) );
  NAND2_X2 U167 ( .A1(StartIn), .A2(n344), .ZN(n398) );
  INV_X4 U168 ( .A(n398), .ZN(n451) );
  XOR2_X2 U169 ( .A(\add/B[9] ), .B(\add/A[9] ), .Z(n348) );
  XOR2_X2 U170 ( .A(n351), .B(n348), .Z(n349) );
  NAND2_X2 U171 ( .A1(StartIn), .A2(n349), .ZN(n397) );
  INV_X4 U172 ( .A(n397), .ZN(n450) );
  NAND2_X2 U173 ( .A1(n351), .A2(n350), .ZN(n353) );
  NAND2_X2 U174 ( .A1(n353), .A2(n352), .ZN(n355) );
  XOR2_X2 U175 ( .A(\add/B[10] ), .B(\add/A[10] ), .Z(n354) );
  XOR2_X2 U176 ( .A(n355), .B(n354), .Z(n356) );
  NAND2_X2 U177 ( .A1(StartIn), .A2(n356), .ZN(n396) );
  INV_X4 U178 ( .A(n396), .ZN(n449) );
  XOR2_X2 U179 ( .A(n386), .B(\add/B[11] ), .Z(n357) );
  XOR2_X2 U180 ( .A(n357), .B(n221), .Z(n358) );
  NAND2_X2 U181 ( .A1(StartIn), .A2(n358), .ZN(n395) );
  INV_X4 U182 ( .A(n395), .ZN(n448) );
  XNOR2_X2 U183 ( .A(\add/B[12] ), .B(\add/A[12] ), .ZN(n360) );
  NAND2_X2 U184 ( .A1(StartIn), .A2(n361), .ZN(n394) );
  INV_X4 U185 ( .A(n394), .ZN(n447) );
  XNOR2_X2 U186 ( .A(\add/B[13] ), .B(\add/A[13] ), .ZN(n363) );
  XNOR2_X2 U187 ( .A(n363), .B(n225), .ZN(n364) );
  NAND2_X2 U188 ( .A1(StartIn), .A2(n364), .ZN(n403) );
  INV_X4 U189 ( .A(n403), .ZN(n446) );
  FA_X1 U190 ( .A(\add/A[14] ), .B(\add/B[14] ), .CI(n227), .S(n365) );
  NAND2_X2 U191 ( .A1(StartIn), .A2(n365), .ZN(n404) );
  INV_X4 U192 ( .A(n404), .ZN(n445) );
  FA_X1 U193 ( .A(\add/A[15] ), .B(\add/B[15] ), .CI(n367), .S(n368) );
  NAND2_X2 U194 ( .A1(StartIn), .A2(n368), .ZN(n393) );
  INV_X4 U195 ( .A(n393), .ZN(n444) );
  FA_X1 U196 ( .A(\add/A[16] ), .B(\add/B[16] ), .CI(n370), .S(n371) );
  NAND2_X2 U197 ( .A1(StartIn), .A2(n371), .ZN(n392) );
  NAND2_X2 U198 ( .A1(n35), .A2(n28), .ZN(n372) );
  NOR4_X2 U199 ( .A1(n372), .A2(\U6/DATA2_5 ), .A3(\U6/DATA2_1 ), .A4(n79), 
        .ZN(n377) );
  NAND4_X2 U200 ( .A1(n32), .A2(n31), .A3(n34), .A4(n33), .ZN(n374) );
  NAND3_X2 U201 ( .A1(n25), .A2(n24), .A3(n26), .ZN(n373) );
  NOR4_X2 U202 ( .A1(n374), .A2(n373), .A3(\U6/DATA2_12 ), .A4(\U6/DATA2_11 ), 
        .ZN(n375) );
  NAND3_X2 U203 ( .A1(n377), .A2(n376), .A3(n375), .ZN(n65) );
  NAND2_X2 U204 ( .A1(StartIn), .A2(n65), .ZN(n437) );
  NAND3_X2 U205 ( .A1(n380), .A2(n379), .A3(n378), .ZN(n383) );
  NAND3_X2 U206 ( .A1(n252), .A2(n245), .A3(n381), .ZN(n382) );
  NOR3_X2 U207 ( .A1(\add/A[18] ), .A2(\add/A[16] ), .A3(\add/A[17] ), .ZN(
        n384) );
  NAND3_X2 U208 ( .A1(n386), .A2(n273), .A3(n385), .ZN(n387) );
  NOR4_X2 U209 ( .A1(n388), .A2(n387), .A3(\add/A[15] ), .A4(\add/A[14] ), 
        .ZN(n389) );
  NAND2_X2 U210 ( .A1(n390), .A2(n389), .ZN(n64) );
  OAI22_X2 U211 ( .A1(n259), .A2(n391), .B1(n24), .B2(n258), .ZN(n84) );
  OAI22_X2 U212 ( .A1(n439), .A2(n392), .B1(n25), .B2(n258), .ZN(n85) );
  OAI22_X2 U213 ( .A1(n259), .A2(n393), .B1(n26), .B2(n437), .ZN(n86) );
  OAI22_X2 U214 ( .A1(n439), .A2(n394), .B1(n29), .B2(n257), .ZN(n89) );
  OAI22_X2 U215 ( .A1(n259), .A2(n395), .B1(n30), .B2(n258), .ZN(n90) );
  OAI22_X2 U216 ( .A1(n439), .A2(n396), .B1(n31), .B2(n437), .ZN(n91) );
  OAI22_X2 U217 ( .A1(n259), .A2(n397), .B1(n32), .B2(n257), .ZN(n92) );
  OAI22_X2 U218 ( .A1(n439), .A2(n398), .B1(n33), .B2(n258), .ZN(n93) );
  OAI22_X2 U219 ( .A1(n259), .A2(n399), .B1(n34), .B2(n437), .ZN(n94) );
  OAI22_X2 U220 ( .A1(n439), .A2(n400), .B1(n40), .B2(n257), .ZN(n100) );
  OAI22_X2 U221 ( .A1(n259), .A2(n401), .B1(n36), .B2(n258), .ZN(n96) );
  OAI22_X2 U222 ( .A1(n439), .A2(n402), .B1(n35), .B2(n437), .ZN(n95) );
  OAI22_X2 U223 ( .A1(n259), .A2(n403), .B1(n28), .B2(n257), .ZN(n88) );
  OAI22_X2 U224 ( .A1(n439), .A2(n404), .B1(n27), .B2(n258), .ZN(n87) );
  INV_X4 U225 ( .A(\add/B[17] ), .ZN(n405) );
  NAND2_X2 U226 ( .A1(n406), .A2(n405), .ZN(n426) );
  INV_X4 U227 ( .A(n426), .ZN(n408) );
  XOR2_X2 U228 ( .A(n423), .B(\add/B[18] ), .Z(n413) );
  NOR3_X2 U229 ( .A1(n408), .A2(n413), .A3(n407), .ZN(n412) );
  NAND2_X2 U230 ( .A1(\add/B[17] ), .A2(\add/A[17] ), .ZN(n427) );
  INV_X4 U231 ( .A(n427), .ZN(n410) );
  INV_X4 U232 ( .A(n413), .ZN(n409) );
  NOR2_X2 U233 ( .A1(n412), .A2(n411), .ZN(n417) );
  NAND2_X2 U234 ( .A1(n408), .A2(n413), .ZN(n416) );
  NOR2_X2 U235 ( .A1(n413), .A2(n427), .ZN(n414) );
  NOR2_X2 U236 ( .A1(n414), .A2(n260), .ZN(n415) );
  NAND3_X2 U237 ( .A1(n417), .A2(n416), .A3(n415), .ZN(n418) );
  INV_X4 U238 ( .A(n418), .ZN(n441) );
  OAI22_X2 U239 ( .A1(n259), .A2(n418), .B1(n23), .B2(n437), .ZN(n83) );
  NAND2_X2 U240 ( .A1(\add/B[18] ), .A2(\add/A[18] ), .ZN(n424) );
  INV_X4 U241 ( .A(n424), .ZN(n421) );
  XOR2_X2 U242 ( .A(n419), .B(\add/B[19] ), .Z(n429) );
  INV_X4 U243 ( .A(n429), .ZN(n420) );
  NAND2_X2 U244 ( .A1(n421), .A2(n420), .ZN(n432) );
  INV_X4 U245 ( .A(\add/B[18] ), .ZN(n422) );
  NAND2_X2 U246 ( .A1(n426), .A2(n425), .ZN(n428) );
  OAI22_X2 U247 ( .A1(n439), .A2(n433), .B1(n21), .B2(n257), .ZN(n82) );
  OAI22_X2 U248 ( .A1(n259), .A2(n434), .B1(n41), .B2(n258), .ZN(n101) );
  OAI22_X2 U249 ( .A1(n439), .A2(n435), .B1(n39), .B2(n437), .ZN(n99) );
  OAI22_X2 U250 ( .A1(n259), .A2(n436), .B1(n38), .B2(n257), .ZN(n98) );
  OAI22_X2 U251 ( .A1(n439), .A2(n438), .B1(n37), .B2(n258), .ZN(n97) );
endmodule


module Cdf_Store ( clock, reset_n, StartIn, ResultIn, StoreAddressIn, WriteBus, 
        WriteAddress, WriteEnable );
  input [19:0] ResultIn;
  input [15:0] StoreAddressIn;
  output [127:0] WriteBus;
  output [15:0] WriteAddress;
  input clock, reset_n, StartIn;
  output WriteEnable;
  wire   \U5/Z_0 , \U5/Z_1 , \U5/Z_2 , \U5/Z_3 , \U5/Z_4 , \U5/Z_5 , \U5/Z_6 ,
         \U5/Z_7 , \U5/Z_8 , \U5/Z_9 , \U5/Z_10 , \U5/Z_11 , \U5/Z_12 ,
         \U5/Z_13 , \U5/Z_14 , \U5/Z_15 , \U5/Z_16 , \U5/Z_17 , \U5/Z_18 ,
         \U5/Z_19 , \U5/DATA1_0 , \U5/DATA1_1 , \U5/DATA1_2 , \U5/DATA1_3 ,
         \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 , \U5/DATA1_7 , \U5/DATA1_8 ,
         \U5/DATA1_9 , \U5/DATA1_10 , \U5/DATA1_11 , \U5/DATA1_12 ,
         \U5/DATA1_13 , \U5/DATA1_14 , \U5/DATA1_15 , \U5/DATA1_16 ,
         \U5/DATA1_17 , \U5/DATA1_18 , \U5/DATA1_19 , \U4/Z_0 , \U4/Z_1 ,
         \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 , \U4/Z_7 , \U4/Z_8 ,
         \U4/Z_9 , \U4/Z_10 , \U4/Z_11 , \U4/Z_12 , \U4/Z_13 , \U4/Z_14 ,
         \U4/Z_15 , \U4/DATA1_0 , \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 ,
         \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 , \U4/DATA1_7 , \U4/DATA1_8 ,
         \U4/DATA1_9 , \U4/DATA1_10 , \U4/DATA1_11 , \U4/DATA1_12 ,
         \U4/DATA1_13 , \U4/DATA1_14 , \U4/DATA1_15 , n443, n444, n445, n446;
  assign \U5/DATA1_0  = ResultIn[0];
  assign \U5/DATA1_1  = ResultIn[1];
  assign \U5/DATA1_2  = ResultIn[2];
  assign \U5/DATA1_3  = ResultIn[3];
  assign \U5/DATA1_4  = ResultIn[4];
  assign \U5/DATA1_5  = ResultIn[5];
  assign \U5/DATA1_6  = ResultIn[6];
  assign \U5/DATA1_7  = ResultIn[7];
  assign \U5/DATA1_8  = ResultIn[8];
  assign \U5/DATA1_9  = ResultIn[9];
  assign \U5/DATA1_10  = ResultIn[10];
  assign \U5/DATA1_11  = ResultIn[11];
  assign \U5/DATA1_12  = ResultIn[12];
  assign \U5/DATA1_13  = ResultIn[13];
  assign \U5/DATA1_14  = ResultIn[14];
  assign \U5/DATA1_15  = ResultIn[15];
  assign \U5/DATA1_16  = ResultIn[16];
  assign \U5/DATA1_17  = ResultIn[17];
  assign \U5/DATA1_18  = ResultIn[18];
  assign \U5/DATA1_19  = ResultIn[19];
  assign \U4/DATA1_0  = StoreAddressIn[0];
  assign \U4/DATA1_1  = StoreAddressIn[1];
  assign \U4/DATA1_2  = StoreAddressIn[2];
  assign \U4/DATA1_3  = StoreAddressIn[3];
  assign \U4/DATA1_4  = StoreAddressIn[4];
  assign \U4/DATA1_5  = StoreAddressIn[5];
  assign \U4/DATA1_6  = StoreAddressIn[6];
  assign \U4/DATA1_7  = StoreAddressIn[7];
  assign \U4/DATA1_8  = StoreAddressIn[8];
  assign \U4/DATA1_9  = StoreAddressIn[9];
  assign \U4/DATA1_10  = StoreAddressIn[10];
  assign \U4/DATA1_11  = StoreAddressIn[11];
  assign \U4/DATA1_12  = StoreAddressIn[12];
  assign \U4/DATA1_13  = StoreAddressIn[13];
  assign \U4/DATA1_14  = StoreAddressIn[14];
  assign \U4/DATA1_15  = StoreAddressIn[15];

  AND2_X1 U131 ( .A1(\U4/DATA1_9 ), .A2(StartIn), .ZN(\U4/Z_9 ) );
  AND2_X1 U132 ( .A1(\U4/DATA1_8 ), .A2(StartIn), .ZN(\U4/Z_8 ) );
  AND2_X1 U133 ( .A1(\U4/DATA1_7 ), .A2(StartIn), .ZN(\U4/Z_7 ) );
  AND2_X1 U134 ( .A1(\U4/DATA1_6 ), .A2(StartIn), .ZN(\U4/Z_6 ) );
  AND2_X1 U135 ( .A1(\U4/DATA1_5 ), .A2(StartIn), .ZN(\U4/Z_5 ) );
  AND2_X1 U136 ( .A1(\U4/DATA1_4 ), .A2(StartIn), .ZN(\U4/Z_4 ) );
  AND2_X1 U137 ( .A1(\U4/DATA1_3 ), .A2(StartIn), .ZN(\U4/Z_3 ) );
  AND2_X1 U138 ( .A1(\U4/DATA1_2 ), .A2(StartIn), .ZN(\U4/Z_2 ) );
  AND2_X1 U139 ( .A1(\U4/DATA1_15 ), .A2(StartIn), .ZN(\U4/Z_15 ) );
  AND2_X1 U140 ( .A1(\U4/DATA1_14 ), .A2(StartIn), .ZN(\U4/Z_14 ) );
  AND2_X1 U141 ( .A1(\U4/DATA1_13 ), .A2(StartIn), .ZN(\U4/Z_13 ) );
  AND2_X1 U142 ( .A1(\U4/DATA1_12 ), .A2(StartIn), .ZN(\U4/Z_12 ) );
  AND2_X1 U143 ( .A1(\U4/DATA1_11 ), .A2(StartIn), .ZN(\U4/Z_11 ) );
  AND2_X1 U144 ( .A1(\U4/DATA1_10 ), .A2(StartIn), .ZN(\U4/Z_10 ) );
  AND2_X1 U145 ( .A1(\U4/DATA1_1 ), .A2(StartIn), .ZN(\U4/Z_1 ) );
  AND2_X1 U146 ( .A1(\U4/DATA1_0 ), .A2(StartIn), .ZN(\U4/Z_0 ) );
  DFFR_X2 WriteEnable_reg ( .D(StartIn), .CK(clock), .RN(n444), .Q(WriteEnable) );
  DFFR_X2 \WriteBus_reg[19]  ( .D(\U5/Z_19 ), .CK(clock), .RN(n444), .Q(
        WriteBus[19]) );
  DFFR_X2 \WriteBus_reg[18]  ( .D(\U5/Z_18 ), .CK(clock), .RN(n444), .Q(
        WriteBus[18]) );
  DFFR_X2 \WriteBus_reg[17]  ( .D(\U5/Z_17 ), .CK(clock), .RN(n444), .Q(
        WriteBus[17]) );
  DFFR_X2 \WriteBus_reg[16]  ( .D(\U5/Z_16 ), .CK(clock), .RN(n444), .Q(
        WriteBus[16]) );
  DFFR_X2 \WriteBus_reg[15]  ( .D(\U5/Z_15 ), .CK(clock), .RN(n444), .Q(
        WriteBus[15]) );
  DFFR_X2 \WriteBus_reg[14]  ( .D(\U5/Z_14 ), .CK(clock), .RN(n444), .Q(
        WriteBus[14]) );
  DFFR_X2 \WriteBus_reg[13]  ( .D(\U5/Z_13 ), .CK(clock), .RN(n444), .Q(
        WriteBus[13]) );
  DFFR_X2 \WriteBus_reg[12]  ( .D(\U5/Z_12 ), .CK(clock), .RN(n444), .Q(
        WriteBus[12]) );
  DFFR_X2 \WriteBus_reg[11]  ( .D(\U5/Z_11 ), .CK(clock), .RN(n443), .Q(
        WriteBus[11]) );
  DFFR_X2 \WriteBus_reg[10]  ( .D(\U5/Z_10 ), .CK(clock), .RN(n443), .Q(
        WriteBus[10]) );
  DFFR_X2 \WriteBus_reg[9]  ( .D(\U5/Z_9 ), .CK(clock), .RN(n443), .Q(
        WriteBus[9]) );
  DFFR_X2 \WriteBus_reg[8]  ( .D(\U5/Z_8 ), .CK(clock), .RN(n443), .Q(
        WriteBus[8]) );
  DFFR_X2 \WriteBus_reg[4]  ( .D(\U5/Z_4 ), .CK(clock), .RN(n443), .Q(
        WriteBus[4]) );
  DFFR_X2 \WriteBus_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .RN(n443), .Q(
        WriteBus[2]) );
  DFFR_X2 \WriteAddress_reg[15]  ( .D(\U4/Z_15 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[15]) );
  DFFR_X2 \WriteAddress_reg[14]  ( .D(\U4/Z_14 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[14]) );
  DFFR_X2 \WriteAddress_reg[13]  ( .D(\U4/Z_13 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[13]) );
  DFFR_X2 \WriteAddress_reg[12]  ( .D(\U4/Z_12 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[12]) );
  DFFR_X2 \WriteAddress_reg[11]  ( .D(\U4/Z_11 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[11]) );
  DFFR_X2 \WriteAddress_reg[10]  ( .D(\U4/Z_10 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[10]) );
  DFFR_X2 \WriteAddress_reg[9]  ( .D(\U4/Z_9 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[9]) );
  DFFR_X2 \WriteAddress_reg[8]  ( .D(\U4/Z_8 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[8]) );
  DFFR_X2 \WriteAddress_reg[7]  ( .D(\U4/Z_7 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[7]) );
  DFFR_X2 \WriteAddress_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[6]) );
  DFFR_X2 \WriteAddress_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[5]) );
  DFFR_X2 \WriteAddress_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[4]) );
  DFFR_X2 \WriteAddress_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[3]) );
  DFFR_X2 \WriteAddress_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[2]) );
  DFFR_X2 \WriteAddress_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[1]) );
  DFFR_X2 \WriteAddress_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[0]) );
  DFFR_X2 \WriteBus_reg[7]  ( .D(\U5/Z_7 ), .CK(clock), .RN(n443), .Q(
        WriteBus[7]) );
  DFFR_X2 \WriteBus_reg[6]  ( .D(\U5/Z_6 ), .CK(clock), .RN(n443), .Q(
        WriteBus[6]) );
  DFFR_X2 \WriteBus_reg[5]  ( .D(\U5/Z_5 ), .CK(clock), .RN(n443), .Q(
        WriteBus[5]) );
  DFFR_X2 \WriteBus_reg[3]  ( .D(\U5/Z_3 ), .CK(clock), .RN(n443), .Q(
        WriteBus[3]) );
  DFFR_X2 \WriteBus_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .RN(n443), .Q(
        WriteBus[1]) );
  DFFR_X2 \WriteBus_reg[0]  ( .D(\U5/Z_0 ), .CK(clock), .RN(n443), .Q(
        WriteBus[0]) );
  INV_X4 U111 ( .A(1'b1), .ZN(WriteBus[20]) );
  INV_X4 U113 ( .A(1'b1), .ZN(WriteBus[21]) );
  INV_X4 U115 ( .A(1'b1), .ZN(WriteBus[22]) );
  INV_X4 U117 ( .A(1'b1), .ZN(WriteBus[23]) );
  INV_X4 U119 ( .A(1'b1), .ZN(WriteBus[24]) );
  INV_X4 U121 ( .A(1'b1), .ZN(WriteBus[25]) );
  INV_X4 U123 ( .A(1'b1), .ZN(WriteBus[26]) );
  INV_X4 U125 ( .A(1'b1), .ZN(WriteBus[27]) );
  INV_X4 U127 ( .A(1'b1), .ZN(WriteBus[28]) );
  INV_X4 U129 ( .A(1'b1), .ZN(WriteBus[29]) );
  INV_X4 U147 ( .A(1'b1), .ZN(WriteBus[30]) );
  INV_X4 U149 ( .A(1'b1), .ZN(WriteBus[31]) );
  INV_X4 U151 ( .A(1'b1), .ZN(WriteBus[32]) );
  INV_X4 U153 ( .A(1'b1), .ZN(WriteBus[33]) );
  INV_X4 U155 ( .A(1'b1), .ZN(WriteBus[34]) );
  INV_X4 U157 ( .A(1'b1), .ZN(WriteBus[35]) );
  INV_X4 U159 ( .A(1'b1), .ZN(WriteBus[36]) );
  INV_X4 U161 ( .A(1'b1), .ZN(WriteBus[37]) );
  INV_X4 U163 ( .A(1'b1), .ZN(WriteBus[38]) );
  INV_X4 U165 ( .A(1'b1), .ZN(WriteBus[39]) );
  INV_X4 U167 ( .A(1'b1), .ZN(WriteBus[40]) );
  INV_X4 U169 ( .A(1'b1), .ZN(WriteBus[41]) );
  INV_X4 U171 ( .A(1'b1), .ZN(WriteBus[42]) );
  INV_X4 U173 ( .A(1'b1), .ZN(WriteBus[43]) );
  INV_X4 U175 ( .A(1'b1), .ZN(WriteBus[44]) );
  INV_X4 U177 ( .A(1'b1), .ZN(WriteBus[45]) );
  INV_X4 U179 ( .A(1'b1), .ZN(WriteBus[46]) );
  INV_X4 U181 ( .A(1'b1), .ZN(WriteBus[47]) );
  INV_X4 U183 ( .A(1'b1), .ZN(WriteBus[48]) );
  INV_X4 U185 ( .A(1'b1), .ZN(WriteBus[49]) );
  INV_X4 U187 ( .A(1'b1), .ZN(WriteBus[50]) );
  INV_X4 U189 ( .A(1'b1), .ZN(WriteBus[51]) );
  INV_X4 U191 ( .A(1'b1), .ZN(WriteBus[52]) );
  INV_X4 U193 ( .A(1'b1), .ZN(WriteBus[53]) );
  INV_X4 U195 ( .A(1'b1), .ZN(WriteBus[54]) );
  INV_X4 U197 ( .A(1'b1), .ZN(WriteBus[55]) );
  INV_X4 U199 ( .A(1'b1), .ZN(WriteBus[56]) );
  INV_X4 U201 ( .A(1'b1), .ZN(WriteBus[57]) );
  INV_X4 U203 ( .A(1'b1), .ZN(WriteBus[58]) );
  INV_X4 U205 ( .A(1'b1), .ZN(WriteBus[59]) );
  INV_X4 U207 ( .A(1'b1), .ZN(WriteBus[60]) );
  INV_X4 U209 ( .A(1'b1), .ZN(WriteBus[61]) );
  INV_X4 U211 ( .A(1'b1), .ZN(WriteBus[62]) );
  INV_X4 U213 ( .A(1'b1), .ZN(WriteBus[63]) );
  INV_X4 U215 ( .A(1'b1), .ZN(WriteBus[64]) );
  INV_X4 U217 ( .A(1'b1), .ZN(WriteBus[65]) );
  INV_X4 U219 ( .A(1'b1), .ZN(WriteBus[66]) );
  INV_X4 U221 ( .A(1'b1), .ZN(WriteBus[67]) );
  INV_X4 U223 ( .A(1'b1), .ZN(WriteBus[68]) );
  INV_X4 U225 ( .A(1'b1), .ZN(WriteBus[69]) );
  INV_X4 U227 ( .A(1'b1), .ZN(WriteBus[70]) );
  INV_X4 U229 ( .A(1'b1), .ZN(WriteBus[71]) );
  INV_X4 U231 ( .A(1'b1), .ZN(WriteBus[72]) );
  INV_X4 U233 ( .A(1'b1), .ZN(WriteBus[73]) );
  INV_X4 U235 ( .A(1'b1), .ZN(WriteBus[74]) );
  INV_X4 U237 ( .A(1'b1), .ZN(WriteBus[75]) );
  INV_X4 U239 ( .A(1'b1), .ZN(WriteBus[76]) );
  INV_X4 U241 ( .A(1'b1), .ZN(WriteBus[77]) );
  INV_X4 U243 ( .A(1'b1), .ZN(WriteBus[78]) );
  INV_X4 U245 ( .A(1'b1), .ZN(WriteBus[79]) );
  INV_X4 U247 ( .A(1'b1), .ZN(WriteBus[80]) );
  INV_X4 U249 ( .A(1'b1), .ZN(WriteBus[81]) );
  INV_X4 U251 ( .A(1'b1), .ZN(WriteBus[82]) );
  INV_X4 U253 ( .A(1'b1), .ZN(WriteBus[83]) );
  INV_X4 U255 ( .A(1'b1), .ZN(WriteBus[84]) );
  INV_X4 U257 ( .A(1'b1), .ZN(WriteBus[85]) );
  INV_X4 U259 ( .A(1'b1), .ZN(WriteBus[86]) );
  INV_X4 U261 ( .A(1'b1), .ZN(WriteBus[87]) );
  INV_X4 U263 ( .A(1'b1), .ZN(WriteBus[88]) );
  INV_X4 U265 ( .A(1'b1), .ZN(WriteBus[89]) );
  INV_X4 U267 ( .A(1'b1), .ZN(WriteBus[90]) );
  INV_X4 U269 ( .A(1'b1), .ZN(WriteBus[91]) );
  INV_X4 U271 ( .A(1'b1), .ZN(WriteBus[92]) );
  INV_X4 U273 ( .A(1'b1), .ZN(WriteBus[93]) );
  INV_X4 U275 ( .A(1'b1), .ZN(WriteBus[94]) );
  INV_X4 U277 ( .A(1'b1), .ZN(WriteBus[95]) );
  INV_X4 U279 ( .A(1'b1), .ZN(WriteBus[96]) );
  INV_X4 U281 ( .A(1'b1), .ZN(WriteBus[97]) );
  INV_X4 U283 ( .A(1'b1), .ZN(WriteBus[98]) );
  INV_X4 U285 ( .A(1'b1), .ZN(WriteBus[99]) );
  INV_X4 U287 ( .A(1'b1), .ZN(WriteBus[100]) );
  INV_X4 U289 ( .A(1'b1), .ZN(WriteBus[101]) );
  INV_X4 U291 ( .A(1'b1), .ZN(WriteBus[102]) );
  INV_X4 U293 ( .A(1'b1), .ZN(WriteBus[103]) );
  INV_X4 U295 ( .A(1'b1), .ZN(WriteBus[104]) );
  INV_X4 U297 ( .A(1'b1), .ZN(WriteBus[105]) );
  INV_X4 U299 ( .A(1'b1), .ZN(WriteBus[106]) );
  INV_X4 U301 ( .A(1'b1), .ZN(WriteBus[107]) );
  INV_X4 U303 ( .A(1'b1), .ZN(WriteBus[108]) );
  INV_X4 U305 ( .A(1'b1), .ZN(WriteBus[109]) );
  INV_X4 U307 ( .A(1'b1), .ZN(WriteBus[110]) );
  INV_X4 U309 ( .A(1'b1), .ZN(WriteBus[111]) );
  INV_X4 U311 ( .A(1'b1), .ZN(WriteBus[112]) );
  INV_X4 U313 ( .A(1'b1), .ZN(WriteBus[113]) );
  INV_X4 U315 ( .A(1'b1), .ZN(WriteBus[114]) );
  INV_X4 U317 ( .A(1'b1), .ZN(WriteBus[115]) );
  INV_X4 U319 ( .A(1'b1), .ZN(WriteBus[116]) );
  INV_X4 U321 ( .A(1'b1), .ZN(WriteBus[117]) );
  INV_X4 U323 ( .A(1'b1), .ZN(WriteBus[118]) );
  INV_X4 U325 ( .A(1'b1), .ZN(WriteBus[119]) );
  INV_X4 U327 ( .A(1'b1), .ZN(WriteBus[120]) );
  INV_X4 U329 ( .A(1'b1), .ZN(WriteBus[121]) );
  INV_X4 U331 ( .A(1'b1), .ZN(WriteBus[122]) );
  INV_X4 U333 ( .A(1'b1), .ZN(WriteBus[123]) );
  INV_X4 U335 ( .A(1'b1), .ZN(WriteBus[124]) );
  INV_X4 U337 ( .A(1'b1), .ZN(WriteBus[125]) );
  INV_X4 U339 ( .A(1'b1), .ZN(WriteBus[126]) );
  INV_X4 U341 ( .A(1'b1), .ZN(WriteBus[127]) );
  INV_X4 U343 ( .A(n446), .ZN(n444) );
  INV_X4 U344 ( .A(n446), .ZN(n443) );
  INV_X4 U345 ( .A(n446), .ZN(n445) );
  INV_X4 U346 ( .A(reset_n), .ZN(n446) );
  AND2_X4 U347 ( .A1(\U5/DATA1_3 ), .A2(StartIn), .ZN(\U5/Z_3 ) );
  AND2_X4 U348 ( .A1(\U5/DATA1_5 ), .A2(StartIn), .ZN(\U5/Z_5 ) );
  AND2_X4 U349 ( .A1(\U5/DATA1_6 ), .A2(StartIn), .ZN(\U5/Z_6 ) );
  AND2_X4 U350 ( .A1(\U5/DATA1_1 ), .A2(StartIn), .ZN(\U5/Z_1 ) );
  AND2_X4 U351 ( .A1(\U5/DATA1_7 ), .A2(StartIn), .ZN(\U5/Z_7 ) );
  AND2_X4 U352 ( .A1(\U5/DATA1_0 ), .A2(StartIn), .ZN(\U5/Z_0 ) );
  AND2_X1 U353 ( .A1(\U5/DATA1_2 ), .A2(StartIn), .ZN(\U5/Z_2 ) );
  AND2_X1 U354 ( .A1(\U5/DATA1_4 ), .A2(StartIn), .ZN(\U5/Z_4 ) );
  AND2_X1 U355 ( .A1(\U5/DATA1_8 ), .A2(StartIn), .ZN(\U5/Z_8 ) );
  AND2_X1 U356 ( .A1(\U5/DATA1_9 ), .A2(StartIn), .ZN(\U5/Z_9 ) );
  AND2_X1 U357 ( .A1(\U5/DATA1_10 ), .A2(StartIn), .ZN(\U5/Z_10 ) );
  AND2_X1 U358 ( .A1(\U5/DATA1_11 ), .A2(StartIn), .ZN(\U5/Z_11 ) );
  AND2_X1 U359 ( .A1(\U5/DATA1_12 ), .A2(StartIn), .ZN(\U5/Z_12 ) );
  AND2_X1 U360 ( .A1(\U5/DATA1_13 ), .A2(StartIn), .ZN(\U5/Z_13 ) );
  AND2_X1 U361 ( .A1(\U5/DATA1_14 ), .A2(StartIn), .ZN(\U5/Z_14 ) );
  AND2_X1 U362 ( .A1(\U5/DATA1_15 ), .A2(StartIn), .ZN(\U5/Z_15 ) );
  AND2_X1 U363 ( .A1(\U5/DATA1_16 ), .A2(StartIn), .ZN(\U5/Z_16 ) );
  AND2_X1 U364 ( .A1(\U5/DATA1_17 ), .A2(StartIn), .ZN(\U5/Z_17 ) );
  AND2_X1 U365 ( .A1(\U5/DATA1_18 ), .A2(StartIn), .ZN(\U5/Z_18 ) );
  AND2_X1 U366 ( .A1(\U5/DATA1_19 ), .A2(StartIn), .ZN(\U5/Z_19 ) );
endmodule


module Cdf_top ( clock, reset_n, start, SP_ReadBus, SP_ReadAddress, 
        WriteEnable, Output_MEMBus, Output_MEMAddress, Cdf_Min, done, 
        input_base_offset, cdf_valid );
  input [127:0] SP_ReadBus;
  output [15:0] SP_ReadAddress;
  output [127:0] Output_MEMBus;
  output [15:0] Output_MEMAddress;
  output [19:0] Cdf_Min;
  input clock, reset_n, start, input_base_offset;
  output WriteEnable, done, cdf_valid;
  wire   n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327,
         start_to_accumlate, start_to_store, n218, n219;
  wire   [19:0] Accumlate;
  wire   [19:0] AccumlateResult;
  wire   [15:0] store_address;
  wire   [15:0] store_address_to_store;

  Cdf_Fetch stage1 ( .clock(clock), .reset_n(n218), .start(start), .ReadBus(
        SP_ReadBus), .ReadAddr(SP_ReadAddress), .AccumlateOut(Accumlate), 
        .StartOut(start_to_accumlate), .StoreAddress(store_address), 
        .input_base_offset(input_base_offset), .done(done) );
  Cdf_Accumlate stage2 ( .clock(clock), .reset_n(n218), .AccumlateIn(Accumlate), .StartIn(start_to_accumlate), .StoreAddressIn(store_address), 
        .AccumlateResult(AccumlateResult), .StoreAddressOut(
        store_address_to_store), .StartOut(start_to_store), .CdfMin(Cdf_Min), 
        .CdfValid(cdf_valid) );
  Cdf_Store stage3 ( .clock(clock), .reset_n(n218), .StartIn(start_to_store), 
        .ResultIn(AccumlateResult), .StoreAddressIn(store_address_to_store), 
        .WriteBus({n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, Output_MEMBus[19:0]}), .WriteAddress(Output_MEMAddress), 
        .WriteEnable(WriteEnable) );
  INV_X4 U1 ( .A(1'b1), .ZN(Output_MEMBus[20]) );
  INV_X4 U3 ( .A(1'b1), .ZN(Output_MEMBus[21]) );
  INV_X4 U5 ( .A(1'b1), .ZN(Output_MEMBus[22]) );
  INV_X4 U7 ( .A(1'b1), .ZN(Output_MEMBus[23]) );
  INV_X4 U9 ( .A(1'b1), .ZN(Output_MEMBus[24]) );
  INV_X4 U11 ( .A(1'b1), .ZN(Output_MEMBus[25]) );
  INV_X4 U13 ( .A(1'b1), .ZN(Output_MEMBus[26]) );
  INV_X4 U15 ( .A(1'b1), .ZN(Output_MEMBus[27]) );
  INV_X4 U17 ( .A(1'b1), .ZN(Output_MEMBus[28]) );
  INV_X4 U19 ( .A(1'b1), .ZN(Output_MEMBus[29]) );
  INV_X4 U21 ( .A(1'b1), .ZN(Output_MEMBus[30]) );
  INV_X4 U23 ( .A(1'b1), .ZN(Output_MEMBus[31]) );
  INV_X4 U25 ( .A(1'b1), .ZN(Output_MEMBus[32]) );
  INV_X4 U27 ( .A(1'b1), .ZN(Output_MEMBus[33]) );
  INV_X4 U29 ( .A(1'b1), .ZN(Output_MEMBus[34]) );
  INV_X4 U31 ( .A(1'b1), .ZN(Output_MEMBus[35]) );
  INV_X4 U33 ( .A(1'b1), .ZN(Output_MEMBus[36]) );
  INV_X4 U35 ( .A(1'b1), .ZN(Output_MEMBus[37]) );
  INV_X4 U37 ( .A(1'b1), .ZN(Output_MEMBus[38]) );
  INV_X4 U39 ( .A(1'b1), .ZN(Output_MEMBus[39]) );
  INV_X4 U41 ( .A(1'b1), .ZN(Output_MEMBus[40]) );
  INV_X4 U43 ( .A(1'b1), .ZN(Output_MEMBus[41]) );
  INV_X4 U45 ( .A(1'b1), .ZN(Output_MEMBus[42]) );
  INV_X4 U47 ( .A(1'b1), .ZN(Output_MEMBus[43]) );
  INV_X4 U49 ( .A(1'b1), .ZN(Output_MEMBus[44]) );
  INV_X4 U51 ( .A(1'b1), .ZN(Output_MEMBus[45]) );
  INV_X4 U53 ( .A(1'b1), .ZN(Output_MEMBus[46]) );
  INV_X4 U55 ( .A(1'b1), .ZN(Output_MEMBus[47]) );
  INV_X4 U57 ( .A(1'b1), .ZN(Output_MEMBus[48]) );
  INV_X4 U59 ( .A(1'b1), .ZN(Output_MEMBus[49]) );
  INV_X4 U61 ( .A(1'b1), .ZN(Output_MEMBus[50]) );
  INV_X4 U63 ( .A(1'b1), .ZN(Output_MEMBus[51]) );
  INV_X4 U65 ( .A(1'b1), .ZN(Output_MEMBus[52]) );
  INV_X4 U67 ( .A(1'b1), .ZN(Output_MEMBus[53]) );
  INV_X4 U69 ( .A(1'b1), .ZN(Output_MEMBus[54]) );
  INV_X4 U71 ( .A(1'b1), .ZN(Output_MEMBus[55]) );
  INV_X4 U73 ( .A(1'b1), .ZN(Output_MEMBus[56]) );
  INV_X4 U75 ( .A(1'b1), .ZN(Output_MEMBus[57]) );
  INV_X4 U77 ( .A(1'b1), .ZN(Output_MEMBus[58]) );
  INV_X4 U79 ( .A(1'b1), .ZN(Output_MEMBus[59]) );
  INV_X4 U81 ( .A(1'b1), .ZN(Output_MEMBus[60]) );
  INV_X4 U83 ( .A(1'b1), .ZN(Output_MEMBus[61]) );
  INV_X4 U85 ( .A(1'b1), .ZN(Output_MEMBus[62]) );
  INV_X4 U87 ( .A(1'b1), .ZN(Output_MEMBus[63]) );
  INV_X4 U89 ( .A(1'b1), .ZN(Output_MEMBus[64]) );
  INV_X4 U91 ( .A(1'b1), .ZN(Output_MEMBus[65]) );
  INV_X4 U93 ( .A(1'b1), .ZN(Output_MEMBus[66]) );
  INV_X4 U95 ( .A(1'b1), .ZN(Output_MEMBus[67]) );
  INV_X4 U97 ( .A(1'b1), .ZN(Output_MEMBus[68]) );
  INV_X4 U99 ( .A(1'b1), .ZN(Output_MEMBus[69]) );
  INV_X4 U101 ( .A(1'b1), .ZN(Output_MEMBus[70]) );
  INV_X4 U103 ( .A(1'b1), .ZN(Output_MEMBus[71]) );
  INV_X4 U105 ( .A(1'b1), .ZN(Output_MEMBus[72]) );
  INV_X4 U107 ( .A(1'b1), .ZN(Output_MEMBus[73]) );
  INV_X4 U109 ( .A(1'b1), .ZN(Output_MEMBus[74]) );
  INV_X4 U111 ( .A(1'b1), .ZN(Output_MEMBus[75]) );
  INV_X4 U113 ( .A(1'b1), .ZN(Output_MEMBus[76]) );
  INV_X4 U115 ( .A(1'b1), .ZN(Output_MEMBus[77]) );
  INV_X4 U117 ( .A(1'b1), .ZN(Output_MEMBus[78]) );
  INV_X4 U119 ( .A(1'b1), .ZN(Output_MEMBus[79]) );
  INV_X4 U121 ( .A(1'b1), .ZN(Output_MEMBus[80]) );
  INV_X4 U123 ( .A(1'b1), .ZN(Output_MEMBus[81]) );
  INV_X4 U125 ( .A(1'b1), .ZN(Output_MEMBus[82]) );
  INV_X4 U127 ( .A(1'b1), .ZN(Output_MEMBus[83]) );
  INV_X4 U129 ( .A(1'b1), .ZN(Output_MEMBus[84]) );
  INV_X4 U131 ( .A(1'b1), .ZN(Output_MEMBus[85]) );
  INV_X4 U133 ( .A(1'b1), .ZN(Output_MEMBus[86]) );
  INV_X4 U135 ( .A(1'b1), .ZN(Output_MEMBus[87]) );
  INV_X4 U137 ( .A(1'b1), .ZN(Output_MEMBus[88]) );
  INV_X4 U139 ( .A(1'b1), .ZN(Output_MEMBus[89]) );
  INV_X4 U141 ( .A(1'b1), .ZN(Output_MEMBus[90]) );
  INV_X4 U143 ( .A(1'b1), .ZN(Output_MEMBus[91]) );
  INV_X4 U145 ( .A(1'b1), .ZN(Output_MEMBus[92]) );
  INV_X4 U147 ( .A(1'b1), .ZN(Output_MEMBus[93]) );
  INV_X4 U149 ( .A(1'b1), .ZN(Output_MEMBus[94]) );
  INV_X4 U151 ( .A(1'b1), .ZN(Output_MEMBus[95]) );
  INV_X4 U153 ( .A(1'b1), .ZN(Output_MEMBus[96]) );
  INV_X4 U155 ( .A(1'b1), .ZN(Output_MEMBus[97]) );
  INV_X4 U157 ( .A(1'b1), .ZN(Output_MEMBus[98]) );
  INV_X4 U159 ( .A(1'b1), .ZN(Output_MEMBus[99]) );
  INV_X4 U161 ( .A(1'b1), .ZN(Output_MEMBus[100]) );
  INV_X4 U163 ( .A(1'b1), .ZN(Output_MEMBus[101]) );
  INV_X4 U165 ( .A(1'b1), .ZN(Output_MEMBus[102]) );
  INV_X4 U167 ( .A(1'b1), .ZN(Output_MEMBus[103]) );
  INV_X4 U169 ( .A(1'b1), .ZN(Output_MEMBus[104]) );
  INV_X4 U171 ( .A(1'b1), .ZN(Output_MEMBus[105]) );
  INV_X4 U173 ( .A(1'b1), .ZN(Output_MEMBus[106]) );
  INV_X4 U175 ( .A(1'b1), .ZN(Output_MEMBus[107]) );
  INV_X4 U177 ( .A(1'b1), .ZN(Output_MEMBus[108]) );
  INV_X4 U179 ( .A(1'b1), .ZN(Output_MEMBus[109]) );
  INV_X4 U181 ( .A(1'b1), .ZN(Output_MEMBus[110]) );
  INV_X4 U183 ( .A(1'b1), .ZN(Output_MEMBus[111]) );
  INV_X4 U185 ( .A(1'b1), .ZN(Output_MEMBus[112]) );
  INV_X4 U187 ( .A(1'b1), .ZN(Output_MEMBus[113]) );
  INV_X4 U189 ( .A(1'b1), .ZN(Output_MEMBus[114]) );
  INV_X4 U191 ( .A(1'b1), .ZN(Output_MEMBus[115]) );
  INV_X4 U193 ( .A(1'b1), .ZN(Output_MEMBus[116]) );
  INV_X4 U195 ( .A(1'b1), .ZN(Output_MEMBus[117]) );
  INV_X4 U197 ( .A(1'b1), .ZN(Output_MEMBus[118]) );
  INV_X4 U199 ( .A(1'b1), .ZN(Output_MEMBus[119]) );
  INV_X4 U201 ( .A(1'b1), .ZN(Output_MEMBus[120]) );
  INV_X4 U203 ( .A(1'b1), .ZN(Output_MEMBus[121]) );
  INV_X4 U205 ( .A(1'b1), .ZN(Output_MEMBus[122]) );
  INV_X4 U207 ( .A(1'b1), .ZN(Output_MEMBus[123]) );
  INV_X4 U209 ( .A(1'b1), .ZN(Output_MEMBus[124]) );
  INV_X4 U211 ( .A(1'b1), .ZN(Output_MEMBus[125]) );
  INV_X4 U213 ( .A(1'b1), .ZN(Output_MEMBus[126]) );
  INV_X4 U215 ( .A(1'b1), .ZN(Output_MEMBus[127]) );
  INV_X4 U217 ( .A(n219), .ZN(n218) );
  INV_X4 U218 ( .A(reset_n), .ZN(n219) );
endmodule


module input_pipeline(
  
);


endmodule


module Output_Fetch_MEM ( clock, reset_n, start, ReadBus, ReadAddress, DataOut, 
        StartOut, StoreAddress, output_base_offset, done );
  input [127:0] ReadBus;
  output [15:0] ReadAddress;
  output [7:0] DataOut;
  output [15:0] StoreAddress;
  input clock, reset_n, start, output_base_offset;
  output StartOut, done;
  wire   n415, n417, n418, n419, n420, n421, n422, n423, n424, U3_U3_Z_0,
         U3_U4_Z_0, U3_U5_Z_0, U3_U5_Z_1, U3_U5_Z_2, U3_U5_Z_3, U6_DATA1_0,
         U6_DATA1_1, U6_DATA1_3, U5_DATA16_0, U5_DATA16_1, U5_DATA16_2,
         U5_DATA16_3, U5_DATA16_4, U5_DATA16_5, U5_DATA16_6, U5_DATA16_7,
         U5_DATA15_0, U5_DATA15_1, U5_DATA15_2, U5_DATA15_3, U5_DATA15_4,
         U5_DATA15_5, U5_DATA15_6, U5_DATA15_7, U5_DATA14_0, U5_DATA14_1,
         U5_DATA14_2, U5_DATA14_3, U5_DATA14_4, U5_DATA14_5, U5_DATA14_6,
         U5_DATA14_7, U5_DATA13_0, U5_DATA13_1, U5_DATA13_2, U5_DATA13_3,
         U5_DATA13_4, U5_DATA13_5, U5_DATA13_6, U5_DATA13_7, U5_DATA12_0,
         U5_DATA12_1, U5_DATA12_2, U5_DATA12_3, U5_DATA12_4, U5_DATA12_5,
         U5_DATA12_6, U5_DATA12_7, U5_DATA11_0, U5_DATA11_1, U5_DATA11_2,
         U5_DATA11_3, U5_DATA11_4, U5_DATA11_5, U5_DATA11_6, U5_DATA11_7,
         U5_DATA10_0, U5_DATA10_1, U5_DATA10_2, U5_DATA10_3, U5_DATA10_4,
         U5_DATA10_5, U5_DATA10_6, U5_DATA10_7, U5_DATA9_0, U5_DATA9_1,
         U5_DATA9_2, U5_DATA9_3, U5_DATA9_4, U5_DATA9_5, U5_DATA9_6,
         U5_DATA9_7, U5_DATA8_0, U5_DATA8_1, U5_DATA8_2, U5_DATA8_3,
         U5_DATA8_4, U5_DATA8_5, U5_DATA8_6, U5_DATA8_7, U5_DATA7_0,
         U5_DATA7_1, U5_DATA7_2, U5_DATA7_3, U5_DATA7_4, U5_DATA7_5,
         U5_DATA7_6, U5_DATA7_7, U5_DATA6_0, U5_DATA6_1, U5_DATA6_2,
         U5_DATA6_3, U5_DATA6_4, U5_DATA6_5, U5_DATA6_6, U5_DATA6_7,
         U5_DATA5_0, U5_DATA5_1, U5_DATA5_2, U5_DATA5_3, U5_DATA5_4,
         U5_DATA5_5, U5_DATA5_6, U5_DATA5_7, U5_DATA4_0, U5_DATA4_1,
         U5_DATA4_2, U5_DATA4_3, U5_DATA4_4, U5_DATA4_5, U5_DATA4_6,
         U5_DATA4_7, U5_DATA3_0, U5_DATA3_1, U5_DATA3_2, U5_DATA3_3,
         U5_DATA3_4, U5_DATA3_5, U5_DATA3_6, U5_DATA3_7, U5_DATA2_0,
         U5_DATA2_1, U5_DATA2_2, U5_DATA2_3, U5_DATA2_4, U5_DATA2_5,
         U5_DATA2_6, U5_DATA2_7, U5_DATA1_0, U5_DATA1_1, U5_DATA1_2,
         U5_DATA1_3, U5_DATA1_4, U5_DATA1_5, U5_DATA1_6, U5_DATA1_7, n147,
         n173, n174, n175, n176, n177, n178, n187, n188, n189, n190, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n268,
         n269, n270, n271, n280, n281, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763;

  DFF_X1 data_in_reg_7_ ( .D(ReadBus[7]), .CK(clock), .Q(U5_DATA1_7) );
  DFF_X1 data_in_reg_6_ ( .D(ReadBus[6]), .CK(clock), .Q(U5_DATA1_6) );
  DFF_X1 data_in_reg_5_ ( .D(ReadBus[5]), .CK(clock), .Q(U5_DATA1_5) );
  DFF_X1 data_in_reg_4_ ( .D(ReadBus[4]), .CK(clock), .Q(U5_DATA1_4) );
  DFF_X1 data_in_reg_3_ ( .D(ReadBus[3]), .CK(clock), .Q(U5_DATA1_3) );
  DFF_X1 data_in_reg_2_ ( .D(ReadBus[2]), .CK(clock), .Q(U5_DATA1_2) );
  DFF_X1 data_in_reg_1_ ( .D(ReadBus[1]), .CK(clock), .Q(U5_DATA1_1) );
  DFF_X1 data_in_reg_0_ ( .D(ReadBus[0]), .CK(clock), .Q(U5_DATA1_0) );
  SDFFR_X2 data_in_reg_107_ ( .D(1'b0), .SI(n642), .SE(ReadBus[107]), .CK(
        clock), .RN(n645), .Q(U5_DATA14_3) );
  SDFFR_X2 data_in_reg_106_ ( .D(1'b0), .SI(n641), .SE(ReadBus[106]), .CK(
        clock), .RN(n645), .Q(U5_DATA14_2) );
  SDFFR_X2 data_in_reg_105_ ( .D(1'b0), .SI(n641), .SE(ReadBus[105]), .CK(
        clock), .RN(n646), .Q(U5_DATA14_1) );
  SDFFR_X2 data_in_reg_104_ ( .D(1'b0), .SI(n642), .SE(ReadBus[104]), .CK(
        clock), .RN(n646), .Q(U5_DATA14_0) );
  SDFFR_X2 data_in_reg_103_ ( .D(1'b0), .SI(n642), .SE(ReadBus[103]), .CK(
        clock), .RN(n646), .Q(U5_DATA13_7) );
  SDFFR_X2 data_in_reg_102_ ( .D(1'b0), .SI(n641), .SE(ReadBus[102]), .CK(
        clock), .RN(n646), .Q(U5_DATA13_6) );
  SDFFR_X2 data_in_reg_101_ ( .D(1'b0), .SI(n641), .SE(ReadBus[101]), .CK(
        clock), .RN(n646), .Q(U5_DATA13_5) );
  SDFFR_X2 data_in_reg_100_ ( .D(1'b0), .SI(n642), .SE(ReadBus[100]), .CK(
        clock), .RN(n646), .Q(U5_DATA13_4) );
  SDFFR_X2 data_in_reg_99_ ( .D(1'b0), .SI(n642), .SE(ReadBus[99]), .CK(clock), 
        .RN(n646), .Q(U5_DATA13_3) );
  SDFFR_X2 data_in_reg_98_ ( .D(1'b0), .SI(n641), .SE(ReadBus[98]), .CK(clock), 
        .RN(n646), .Q(U5_DATA13_2) );
  SDFFR_X2 data_in_reg_17_ ( .D(1'b0), .SI(n641), .SE(ReadBus[17]), .CK(clock), 
        .RN(n646), .Q(U5_DATA3_1) );
  SDFFR_X2 data_in_reg_97_ ( .D(1'b0), .SI(n642), .SE(ReadBus[97]), .CK(clock), 
        .RN(n646), .Q(U5_DATA13_1) );
  SDFFR_X2 data_in_reg_96_ ( .D(1'b0), .SI(n642), .SE(ReadBus[96]), .CK(clock), 
        .RN(n646), .Q(U5_DATA13_0) );
  SDFFR_X2 data_in_reg_95_ ( .D(1'b0), .SI(n641), .SE(ReadBus[95]), .CK(clock), 
        .RN(n646), .Q(U5_DATA12_7) );
  SDFFR_X2 data_in_reg_94_ ( .D(1'b0), .SI(n641), .SE(ReadBus[94]), .CK(clock), 
        .RN(n646), .Q(U5_DATA12_6) );
  SDFFR_X2 data_in_reg_93_ ( .D(1'b0), .SI(n642), .SE(ReadBus[93]), .CK(clock), 
        .RN(n646), .Q(U5_DATA12_5) );
  SDFFR_X2 data_in_reg_92_ ( .D(1'b0), .SI(n642), .SE(ReadBus[92]), .CK(clock), 
        .RN(n646), .Q(U5_DATA12_4) );
  SDFFR_X2 data_in_reg_91_ ( .D(1'b0), .SI(n641), .SE(ReadBus[91]), .CK(clock), 
        .RN(n646), .Q(U5_DATA12_3) );
  SDFFR_X2 data_in_reg_90_ ( .D(1'b0), .SI(n641), .SE(ReadBus[90]), .CK(clock), 
        .RN(n646), .Q(U5_DATA12_2) );
  SDFFR_X2 data_in_reg_89_ ( .D(1'b0), .SI(n642), .SE(ReadBus[89]), .CK(clock), 
        .RN(n646), .Q(U5_DATA12_1) );
  SDFFR_X2 data_in_reg_88_ ( .D(1'b0), .SI(n642), .SE(ReadBus[88]), .CK(clock), 
        .RN(n646), .Q(U5_DATA12_0) );
  SDFFR_X2 data_in_reg_16_ ( .D(1'b0), .SI(n641), .SE(ReadBus[16]), .CK(clock), 
        .RN(n646), .Q(U5_DATA3_0) );
  SDFFR_X2 data_in_reg_87_ ( .D(1'b0), .SI(n642), .SE(ReadBus[87]), .CK(clock), 
        .RN(n646), .Q(U5_DATA11_7) );
  SDFFR_X2 data_in_reg_86_ ( .D(1'b0), .SI(n641), .SE(ReadBus[86]), .CK(clock), 
        .RN(n646), .Q(U5_DATA11_6) );
  SDFFR_X2 data_in_reg_85_ ( .D(1'b0), .SI(n642), .SE(ReadBus[85]), .CK(clock), 
        .RN(n646), .Q(U5_DATA11_5) );
  SDFFR_X2 data_in_reg_84_ ( .D(1'b0), .SI(n641), .SE(ReadBus[84]), .CK(clock), 
        .RN(n646), .Q(U5_DATA11_4) );
  SDFFR_X2 data_in_reg_83_ ( .D(1'b0), .SI(n642), .SE(ReadBus[83]), .CK(clock), 
        .RN(n646), .Q(U5_DATA11_3) );
  SDFFR_X2 data_in_reg_82_ ( .D(1'b0), .SI(n641), .SE(ReadBus[82]), .CK(clock), 
        .RN(n646), .Q(U5_DATA11_2) );
  SDFFR_X2 data_in_reg_81_ ( .D(1'b0), .SI(n642), .SE(ReadBus[81]), .CK(clock), 
        .RN(n646), .Q(U5_DATA11_1) );
  SDFFR_X2 data_in_reg_80_ ( .D(1'b0), .SI(n641), .SE(ReadBus[80]), .CK(clock), 
        .RN(n646), .Q(U5_DATA11_0) );
  SDFFR_X2 data_in_reg_79_ ( .D(1'b0), .SI(n642), .SE(ReadBus[79]), .CK(clock), 
        .RN(n646), .Q(U5_DATA10_7) );
  SDFFR_X2 data_in_reg_78_ ( .D(1'b0), .SI(n641), .SE(ReadBus[78]), .CK(clock), 
        .RN(n647), .Q(U5_DATA10_6) );
  SDFFR_X2 data_in_reg_15_ ( .D(1'b0), .SI(n642), .SE(ReadBus[15]), .CK(clock), 
        .RN(n647), .Q(U5_DATA2_7) );
  SDFFR_X2 data_in_reg_77_ ( .D(1'b0), .SI(n641), .SE(ReadBus[77]), .CK(clock), 
        .RN(n647), .Q(U5_DATA10_5) );
  SDFFR_X2 data_in_reg_76_ ( .D(1'b0), .SI(n642), .SE(ReadBus[76]), .CK(clock), 
        .RN(n647), .Q(U5_DATA10_4) );
  SDFFR_X2 data_in_reg_75_ ( .D(1'b0), .SI(n641), .SE(ReadBus[75]), .CK(clock), 
        .RN(n647), .Q(U5_DATA10_3) );
  SDFFR_X2 data_in_reg_74_ ( .D(1'b0), .SI(n642), .SE(ReadBus[74]), .CK(clock), 
        .RN(n647), .Q(U5_DATA10_2) );
  SDFFR_X2 data_in_reg_73_ ( .D(1'b0), .SI(n641), .SE(ReadBus[73]), .CK(clock), 
        .RN(n647), .Q(U5_DATA10_1) );
  SDFFR_X2 data_in_reg_72_ ( .D(1'b0), .SI(n642), .SE(ReadBus[72]), .CK(clock), 
        .RN(n647), .Q(U5_DATA10_0) );
  SDFFR_X2 data_in_reg_71_ ( .D(1'b0), .SI(n641), .SE(ReadBus[71]), .CK(clock), 
        .RN(n647), .Q(U5_DATA9_7) );
  SDFFR_X2 data_in_reg_70_ ( .D(1'b0), .SI(n642), .SE(ReadBus[70]), .CK(clock), 
        .RN(n647), .Q(U5_DATA9_6) );
  SDFFR_X2 data_in_reg_69_ ( .D(1'b0), .SI(n641), .SE(ReadBus[69]), .CK(clock), 
        .RN(n647), .Q(U5_DATA9_5) );
  SDFFR_X2 data_in_reg_68_ ( .D(1'b0), .SI(n642), .SE(ReadBus[68]), .CK(clock), 
        .RN(n647), .Q(U5_DATA9_4) );
  SDFFR_X2 data_in_reg_14_ ( .D(1'b0), .SI(n641), .SE(ReadBus[14]), .CK(clock), 
        .RN(n647), .Q(U5_DATA2_6) );
  SDFFR_X2 data_in_reg_67_ ( .D(1'b0), .SI(n641), .SE(ReadBus[67]), .CK(clock), 
        .RN(n647), .Q(U5_DATA9_3) );
  SDFFR_X2 data_in_reg_66_ ( .D(1'b0), .SI(n642), .SE(ReadBus[66]), .CK(clock), 
        .RN(n647), .Q(U5_DATA9_2) );
  SDFFR_X2 data_in_reg_65_ ( .D(1'b0), .SI(n642), .SE(ReadBus[65]), .CK(clock), 
        .RN(n647), .Q(U5_DATA9_1) );
  SDFFR_X2 data_in_reg_64_ ( .D(1'b0), .SI(n641), .SE(ReadBus[64]), .CK(clock), 
        .RN(n647), .Q(U5_DATA9_0) );
  SDFFR_X2 data_in_reg_63_ ( .D(1'b0), .SI(n642), .SE(ReadBus[63]), .CK(clock), 
        .RN(n647), .Q(U5_DATA8_7) );
  SDFFR_X2 data_in_reg_62_ ( .D(1'b0), .SI(n641), .SE(ReadBus[62]), .CK(clock), 
        .RN(n647), .Q(U5_DATA8_6) );
  SDFFR_X2 data_in_reg_61_ ( .D(1'b0), .SI(n641), .SE(ReadBus[61]), .CK(clock), 
        .RN(n647), .Q(U5_DATA8_5) );
  SDFFR_X2 data_in_reg_60_ ( .D(1'b0), .SI(n642), .SE(ReadBus[60]), .CK(clock), 
        .RN(n647), .Q(U5_DATA8_4) );
  SDFFR_X2 data_in_reg_59_ ( .D(1'b0), .SI(n642), .SE(ReadBus[59]), .CK(clock), 
        .RN(n647), .Q(U5_DATA8_3) );
  SDFFR_X2 data_in_reg_58_ ( .D(1'b0), .SI(n641), .SE(ReadBus[58]), .CK(clock), 
        .RN(n647), .Q(U5_DATA8_2) );
  SDFFR_X2 data_in_reg_13_ ( .D(1'b0), .SI(n641), .SE(ReadBus[13]), .CK(clock), 
        .RN(n647), .Q(U5_DATA2_5) );
  SDFFR_X2 data_in_reg_57_ ( .D(1'b0), .SI(n642), .SE(ReadBus[57]), .CK(clock), 
        .RN(n647), .Q(U5_DATA8_1) );
  SDFFR_X2 data_in_reg_56_ ( .D(1'b0), .SI(n641), .SE(ReadBus[56]), .CK(clock), 
        .RN(n647), .Q(U5_DATA8_0) );
  SDFFR_X2 data_in_reg_55_ ( .D(1'b0), .SI(n642), .SE(ReadBus[55]), .CK(clock), 
        .RN(n647), .Q(U5_DATA7_7) );
  SDFFR_X2 data_in_reg_54_ ( .D(1'b0), .SI(n642), .SE(ReadBus[54]), .CK(clock), 
        .RN(n647), .Q(U5_DATA7_6) );
  SDFFR_X2 data_in_reg_53_ ( .D(1'b0), .SI(n641), .SE(ReadBus[53]), .CK(clock), 
        .RN(n648), .Q(U5_DATA7_5) );
  SDFFR_X2 data_in_reg_52_ ( .D(1'b0), .SI(n642), .SE(ReadBus[52]), .CK(clock), 
        .RN(n648), .Q(U5_DATA7_4) );
  SDFFR_X2 data_in_reg_51_ ( .D(1'b0), .SI(n641), .SE(ReadBus[51]), .CK(clock), 
        .RN(n648), .Q(U5_DATA7_3) );
  SDFFR_X2 data_in_reg_50_ ( .D(1'b0), .SI(n642), .SE(ReadBus[50]), .CK(clock), 
        .RN(n648), .Q(U5_DATA7_2) );
  SDFFR_X2 data_in_reg_49_ ( .D(1'b0), .SI(n641), .SE(ReadBus[49]), .CK(clock), 
        .RN(n648), .Q(U5_DATA7_1) );
  SDFFR_X2 data_in_reg_48_ ( .D(1'b0), .SI(n641), .SE(ReadBus[48]), .CK(clock), 
        .RN(n648), .Q(U5_DATA7_0) );
  SDFFR_X2 data_in_reg_12_ ( .D(1'b0), .SI(n642), .SE(ReadBus[12]), .CK(clock), 
        .RN(n648), .Q(U5_DATA2_4) );
  SDFFR_X2 data_in_reg_47_ ( .D(1'b0), .SI(n642), .SE(ReadBus[47]), .CK(clock), 
        .RN(n648), .Q(U5_DATA6_7) );
  SDFFR_X2 data_in_reg_46_ ( .D(1'b0), .SI(n641), .SE(ReadBus[46]), .CK(clock), 
        .RN(n648), .Q(U5_DATA6_6) );
  SDFFR_X2 data_in_reg_45_ ( .D(1'b0), .SI(n641), .SE(ReadBus[45]), .CK(clock), 
        .RN(n648), .Q(U5_DATA6_5) );
  SDFFR_X2 data_in_reg_44_ ( .D(1'b0), .SI(n642), .SE(ReadBus[44]), .CK(clock), 
        .RN(n648), .Q(U5_DATA6_4) );
  SDFFR_X2 data_in_reg_43_ ( .D(1'b0), .SI(n642), .SE(ReadBus[43]), .CK(clock), 
        .RN(n648), .Q(U5_DATA6_3) );
  SDFFR_X2 data_in_reg_42_ ( .D(1'b0), .SI(n641), .SE(ReadBus[42]), .CK(clock), 
        .RN(n648), .Q(U5_DATA6_2) );
  SDFFR_X2 data_in_reg_41_ ( .D(1'b0), .SI(n641), .SE(ReadBus[41]), .CK(clock), 
        .RN(n648), .Q(U5_DATA6_1) );
  SDFFR_X2 data_in_reg_40_ ( .D(1'b0), .SI(n642), .SE(ReadBus[40]), .CK(clock), 
        .RN(n648), .Q(U5_DATA6_0) );
  SDFFR_X2 data_in_reg_39_ ( .D(1'b0), .SI(n642), .SE(ReadBus[39]), .CK(clock), 
        .RN(n648), .Q(U5_DATA5_7) );
  SDFFR_X2 data_in_reg_38_ ( .D(1'b0), .SI(n641), .SE(ReadBus[38]), .CK(clock), 
        .RN(n648), .Q(U5_DATA5_6) );
  SDFFR_X2 data_in_reg_11_ ( .D(1'b0), .SI(n641), .SE(ReadBus[11]), .CK(clock), 
        .RN(n648), .Q(U5_DATA2_3) );
  SDFFR_X2 data_in_reg_37_ ( .D(1'b0), .SI(n642), .SE(ReadBus[37]), .CK(clock), 
        .RN(n648), .Q(U5_DATA5_5) );
  SDFFR_X2 data_in_reg_36_ ( .D(1'b0), .SI(n642), .SE(ReadBus[36]), .CK(clock), 
        .RN(n648), .Q(U5_DATA5_4) );
  SDFFR_X2 data_in_reg_35_ ( .D(1'b0), .SI(n641), .SE(ReadBus[35]), .CK(clock), 
        .RN(n648), .Q(U5_DATA5_3) );
  SDFFR_X2 data_in_reg_34_ ( .D(1'b0), .SI(n642), .SE(ReadBus[34]), .CK(clock), 
        .RN(n648), .Q(U5_DATA5_2) );
  SDFFR_X2 data_in_reg_33_ ( .D(1'b0), .SI(n641), .SE(ReadBus[33]), .CK(clock), 
        .RN(n647), .Q(U5_DATA5_1) );
  SDFFR_X2 data_in_reg_32_ ( .D(1'b0), .SI(n641), .SE(ReadBus[32]), .CK(clock), 
        .RN(n648), .Q(U5_DATA5_0) );
  SDFFR_X2 data_in_reg_31_ ( .D(1'b0), .SI(n642), .SE(ReadBus[31]), .CK(clock), 
        .RN(n648), .Q(U5_DATA4_7) );
  SDFFR_X2 data_in_reg_30_ ( .D(1'b0), .SI(n642), .SE(ReadBus[30]), .CK(clock), 
        .RN(n648), .Q(U5_DATA4_6) );
  SDFFR_X2 data_in_reg_29_ ( .D(1'b0), .SI(n641), .SE(ReadBus[29]), .CK(clock), 
        .RN(n648), .Q(U5_DATA4_5) );
  SDFFR_X2 data_in_reg_28_ ( .D(1'b0), .SI(n641), .SE(ReadBus[28]), .CK(clock), 
        .RN(n648), .Q(U5_DATA4_4) );
  SDFFR_X2 data_in_reg_10_ ( .D(1'b0), .SI(n642), .SE(ReadBus[10]), .CK(clock), 
        .RN(n648), .Q(U5_DATA2_2) );
  SDFFR_X2 data_in_reg_27_ ( .D(1'b0), .SI(n642), .SE(ReadBus[27]), .CK(clock), 
        .RN(n648), .Q(U5_DATA4_3) );
  SDFFR_X2 data_in_reg_26_ ( .D(1'b0), .SI(n641), .SE(ReadBus[26]), .CK(clock), 
        .RN(n649), .Q(U5_DATA4_2) );
  SDFFR_X2 data_in_reg_25_ ( .D(1'b0), .SI(n642), .SE(ReadBus[25]), .CK(clock), 
        .RN(n649), .Q(U5_DATA4_1) );
  SDFFR_X2 data_in_reg_24_ ( .D(1'b0), .SI(n641), .SE(ReadBus[24]), .CK(clock), 
        .RN(n649), .Q(U5_DATA4_0) );
  SDFFR_X2 data_in_reg_23_ ( .D(1'b0), .SI(n642), .SE(ReadBus[23]), .CK(clock), 
        .RN(n649), .Q(U5_DATA3_7) );
  SDFFR_X2 data_in_reg_22_ ( .D(1'b0), .SI(n641), .SE(ReadBus[22]), .CK(clock), 
        .RN(n649), .Q(U5_DATA3_6) );
  SDFFR_X2 data_in_reg_21_ ( .D(1'b0), .SI(n642), .SE(ReadBus[21]), .CK(clock), 
        .RN(n649), .Q(U5_DATA3_5) );
  SDFFR_X2 data_in_reg_20_ ( .D(1'b0), .SI(n641), .SE(ReadBus[20]), .CK(clock), 
        .RN(n649), .Q(U5_DATA3_4) );
  SDFFR_X2 data_in_reg_127_ ( .D(1'b0), .SI(n642), .SE(ReadBus[127]), .CK(
        clock), .RN(n649), .Q(U5_DATA16_7) );
  SDFFR_X2 data_in_reg_126_ ( .D(1'b0), .SI(n641), .SE(ReadBus[126]), .CK(
        clock), .RN(n649), .Q(U5_DATA16_6) );
  SDFFR_X2 data_in_reg_125_ ( .D(1'b0), .SI(n642), .SE(ReadBus[125]), .CK(
        clock), .RN(n649), .Q(U5_DATA16_5) );
  SDFFR_X2 data_in_reg_124_ ( .D(1'b0), .SI(n641), .SE(ReadBus[124]), .CK(
        clock), .RN(n649), .Q(U5_DATA16_4) );
  SDFFR_X2 data_in_reg_123_ ( .D(1'b0), .SI(n642), .SE(ReadBus[123]), .CK(
        clock), .RN(n649), .Q(U5_DATA16_3) );
  SDFFR_X2 data_in_reg_122_ ( .D(1'b0), .SI(n641), .SE(ReadBus[122]), .CK(
        clock), .RN(n649), .Q(U5_DATA16_2) );
  SDFFR_X2 data_in_reg_121_ ( .D(1'b0), .SI(n642), .SE(ReadBus[121]), .CK(
        clock), .RN(n649), .Q(U5_DATA16_1) );
  SDFFR_X2 data_in_reg_120_ ( .D(1'b0), .SI(n641), .SE(ReadBus[120]), .CK(
        clock), .RN(n649), .Q(U5_DATA16_0) );
  SDFFR_X2 data_in_reg_119_ ( .D(1'b0), .SI(n641), .SE(ReadBus[119]), .CK(
        clock), .RN(n649), .Q(U5_DATA15_7) );
  SDFFR_X2 data_in_reg_118_ ( .D(1'b0), .SI(n642), .SE(ReadBus[118]), .CK(
        clock), .RN(n649), .Q(U5_DATA15_6) );
  SDFFR_X2 data_in_reg_19_ ( .D(1'b0), .SI(n641), .SE(ReadBus[19]), .CK(clock), 
        .RN(n649), .Q(U5_DATA3_3) );
  SDFFR_X2 data_in_reg_117_ ( .D(1'b0), .SI(n642), .SE(ReadBus[117]), .CK(
        clock), .RN(n649), .Q(U5_DATA15_5) );
  SDFFR_X2 data_in_reg_116_ ( .D(1'b0), .SI(n641), .SE(ReadBus[116]), .CK(
        clock), .RN(n649), .Q(U5_DATA15_4) );
  SDFFR_X2 data_in_reg_115_ ( .D(1'b0), .SI(n642), .SE(ReadBus[115]), .CK(
        clock), .RN(n649), .Q(U5_DATA15_3) );
  SDFFR_X2 data_in_reg_114_ ( .D(1'b0), .SI(n642), .SE(ReadBus[114]), .CK(
        clock), .RN(n649), .Q(U5_DATA15_2) );
  SDFFR_X2 data_in_reg_113_ ( .D(1'b0), .SI(n641), .SE(ReadBus[113]), .CK(
        clock), .RN(n649), .Q(U5_DATA15_1) );
  SDFFR_X2 data_in_reg_112_ ( .D(1'b0), .SI(n642), .SE(ReadBus[112]), .CK(
        clock), .RN(n649), .Q(U5_DATA15_0) );
  SDFFR_X2 data_in_reg_111_ ( .D(1'b0), .SI(n641), .SE(ReadBus[111]), .CK(
        clock), .RN(n649), .Q(U5_DATA14_7) );
  SDFFR_X2 data_in_reg_110_ ( .D(1'b0), .SI(n642), .SE(ReadBus[110]), .CK(
        clock), .RN(n649), .Q(U5_DATA14_6) );
  SDFFR_X2 data_in_reg_109_ ( .D(1'b0), .SI(n641), .SE(ReadBus[109]), .CK(
        clock), .RN(n649), .Q(U5_DATA14_5) );
  SDFFR_X2 data_in_reg_108_ ( .D(1'b0), .SI(n642), .SE(ReadBus[108]), .CK(
        clock), .RN(n649), .Q(U5_DATA14_4) );
  SDFFR_X2 data_in_reg_18_ ( .D(1'b0), .SI(n641), .SE(ReadBus[18]), .CK(clock), 
        .RN(n649), .Q(U5_DATA3_2) );
  SDFFR_X2 data_in_reg_9_ ( .D(1'b0), .SI(start), .SE(ReadBus[9]), .CK(clock), 
        .RN(reset_n), .Q(U5_DATA2_1) );
  SDFFR_X2 data_in_reg_8_ ( .D(1'b0), .SI(start), .SE(ReadBus[8]), .CK(clock), 
        .RN(n645), .Q(U5_DATA2_0) );
  NAND4_X2 U143 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(n174) );
  NAND4_X2 U148 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(n173) );
  NAND4_X2 U153 ( .A1(n201), .A2(n202), .A3(n203), .A4(n204), .ZN(n200) );
  NAND4_X2 U158 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(n199) );
  NAND4_X2 U163 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(n210) );
  NAND4_X2 U168 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(n209) );
  NAND4_X2 U173 ( .A1(n221), .A2(n222), .A3(n223), .A4(n224), .ZN(n220) );
  NAND4_X2 U178 ( .A1(n225), .A2(n226), .A3(n227), .A4(n228), .ZN(n219) );
  NAND4_X2 U183 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(n230) );
  NAND4_X2 U188 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(n229) );
  NAND4_X2 U193 ( .A1(n241), .A2(n242), .A3(n243), .A4(n244), .ZN(n240) );
  NAND4_X2 U198 ( .A1(n245), .A2(n246), .A3(n247), .A4(n248), .ZN(n239) );
  NAND4_X2 U203 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(n250) );
  NAND4_X2 U208 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(n249) );
  NAND4_X2 U213 ( .A1(n261), .A2(n262), .A3(n263), .A4(n264), .ZN(n260) );
  NAND4_X2 U225 ( .A1(n268), .A2(n269), .A3(n270), .A4(n271), .ZN(n259) );
  OR2_X1 U284 ( .A1(n173), .A2(n174), .ZN(DataOut[7]) );
  OR2_X1 U285 ( .A1(n199), .A2(n200), .ZN(DataOut[6]) );
  OR2_X1 U286 ( .A1(n209), .A2(n210), .ZN(DataOut[5]) );
  OR2_X1 U287 ( .A1(n219), .A2(n220), .ZN(DataOut[4]) );
  OR2_X1 U288 ( .A1(n229), .A2(n230), .ZN(DataOut[3]) );
  OR2_X1 U289 ( .A1(n239), .A2(n240), .ZN(DataOut[2]) );
  OR2_X1 U290 ( .A1(n249), .A2(n250), .ZN(DataOut[1]) );
  OR2_X1 U291 ( .A1(n259), .A2(n260), .ZN(DataOut[0]) );
  DFFR_X2 ReadAddress_reg_2_ ( .D(n762), .CK(clock), .RN(reset_n), .Q(
        ReadAddress[2]), .QN(n629) );
  DFFR_X2 done8_reg ( .D(n417), .CK(clock), .RN(n644), .Q(n415) );
  DFFR_X2 done7_reg ( .D(n418), .CK(clock), .RN(reset_n), .Q(n417) );
  DFFR_X2 done6_reg ( .D(n419), .CK(clock), .RN(reset_n), .Q(n418) );
  DFFR_X2 done5_reg ( .D(n420), .CK(clock), .RN(n645), .Q(n419) );
  DFFR_X2 done4_reg ( .D(n421), .CK(clock), .RN(n645), .Q(n420) );
  DFFR_X2 done3_reg ( .D(n422), .CK(clock), .RN(n648), .Q(n421) );
  DFFR_X2 done2_reg ( .D(n423), .CK(clock), .RN(n649), .Q(n422) );
  DFFR_X2 done1_reg ( .D(n424), .CK(clock), .RN(n648), .Q(n423) );
  DFFR_X2 StoreAddress_reg_15_ ( .D(ReadAddress[15]), .CK(clock), .RN(n649), 
        .Q(StoreAddress[15]) );
  DFFR_X2 StoreAddress_reg_2_ ( .D(ReadAddress[2]), .CK(clock), .RN(reset_n), 
        .Q(StoreAddress[2]) );
  DFFR_X2 StoreAddress_reg_6_ ( .D(ReadAddress[6]), .CK(clock), .RN(n644), .Q(
        StoreAddress[6]) );
  DFFR_X2 StoreAddress_reg_4_ ( .D(ReadAddress[4]), .CK(clock), .RN(n644), .Q(
        StoreAddress[4]) );
  DFFR_X2 StoreAddress_reg_0_ ( .D(ReadAddress[0]), .CK(clock), .RN(n646), .Q(
        StoreAddress[0]) );
  DFFR_X2 StoreAddress_reg_12_ ( .D(ReadAddress[12]), .CK(clock), .RN(n645), 
        .Q(StoreAddress[12]) );
  DFFR_X2 StoreAddress_reg_8_ ( .D(ReadAddress[8]), .CK(clock), .RN(n644), .Q(
        StoreAddress[8]) );
  DFFR_X2 StoreAddress_reg_1_ ( .D(ReadAddress[1]), .CK(clock), .RN(reset_n), 
        .Q(StoreAddress[1]) );
  DFFR_X2 StoreAddress_reg_5_ ( .D(ReadAddress[5]), .CK(clock), .RN(n644), .Q(
        StoreAddress[5]) );
  DFFR_X2 StoreAddress_reg_3_ ( .D(ReadAddress[3]), .CK(clock), .RN(reset_n), 
        .Q(StoreAddress[3]) );
  DFFR_X2 StoreAddress_reg_10_ ( .D(ReadAddress[10]), .CK(clock), .RN(n645), 
        .Q(StoreAddress[10]) );
  DFFR_X2 StoreAddress_reg_14_ ( .D(ReadAddress[14]), .CK(clock), .RN(n645), 
        .Q(StoreAddress[14]) );
  DFFR_X2 StoreAddress_reg_13_ ( .D(ReadAddress[13]), .CK(clock), .RN(n645), 
        .Q(StoreAddress[13]) );
  DFFR_X2 StoreAddress_reg_11_ ( .D(ReadAddress[11]), .CK(clock), .RN(n645), 
        .Q(StoreAddress[11]) );
  DFFR_X2 StoreAddress_reg_7_ ( .D(ReadAddress[7]), .CK(clock), .RN(n644), .Q(
        StoreAddress[7]) );
  DFFR_X2 StoreAddress_reg_9_ ( .D(ReadAddress[9]), .CK(clock), .RN(n644), .Q(
        StoreAddress[9]) );
  DFFR_X2 StartOut_reg ( .D(U3_U3_Z_0), .CK(clock), .RN(n645), .Q(StartOut) );
  DFFR_X2 done0_reg ( .D(U3_U4_Z_0), .CK(clock), .RN(n644), .Q(n424) );
  DFFR_X2 short_count_reg_0_ ( .D(U3_U5_Z_0), .CK(clock), .RN(reset_n), .Q(
        U6_DATA1_0), .QN(n742) );
  DFFR_X2 short_count_reg_1_ ( .D(U3_U5_Z_1), .CK(clock), .RN(reset_n), .Q(
        U6_DATA1_1), .QN(n739) );
  DFFR_X2 done_reg ( .D(n415), .CK(clock), .RN(reset_n), .Q(done) );
  DFFR_X2 ReadAddress_reg_6_ ( .D(n758), .CK(clock), .RN(n644), .Q(
        ReadAddress[6]), .QN(n682) );
  DFFR_X2 ReadAddress_reg_8_ ( .D(n756), .CK(clock), .RN(n644), .Q(
        ReadAddress[8]), .QN(n714) );
  DFFR_X2 ReadAddress_reg_14_ ( .D(n750), .CK(clock), .RN(n645), .Q(
        ReadAddress[14]), .QN(n727) );
  DFFR_X2 ReadAddress_reg_4_ ( .D(n760), .CK(clock), .RN(reset_n), .Q(
        ReadAddress[4]), .QN(n673) );
  DFFR_X2 ReadAddress_reg_10_ ( .D(n754), .CK(clock), .RN(n644), .Q(
        ReadAddress[10]), .QN(n713) );
  DFFR_X2 ReadAddress_reg_12_ ( .D(n752), .CK(clock), .RN(n645), .Q(
        ReadAddress[12]), .QN(n705) );
  DFFR_X2 short_count_reg_3_ ( .D(U3_U5_Z_3), .CK(clock), .RN(reset_n), .Q(
        U6_DATA1_3), .QN(n744) );
  DFFR_X2 short_count_reg_2_ ( .D(U3_U5_Z_2), .CK(clock), .RN(reset_n), .Q(
        n741), .QN(n746) );
  DFFR_X2 ReadAddress_reg_15_ ( .D(n280), .CK(clock), .RN(reset_n), .Q(
        ReadAddress[15]), .QN(n147) );
  DFFR_X2 ReadAddress_reg_0_ ( .D(n281), .CK(clock), .RN(n645), .Q(
        ReadAddress[0]), .QN(n660) );
  DFFR_X2 ReadAddress_reg_13_ ( .D(n751), .CK(clock), .RN(n645), .Q(
        ReadAddress[13]), .QN(n711) );
  DFFR_X2 ReadAddress_reg_11_ ( .D(n753), .CK(clock), .RN(n645), .Q(
        ReadAddress[11]), .QN(n653) );
  DFFR_X2 ReadAddress_reg_9_ ( .D(n755), .CK(clock), .RN(n644), .Q(
        ReadAddress[9]), .QN(n652) );
  DFFR_X2 ReadAddress_reg_7_ ( .D(n757), .CK(clock), .RN(n644), .Q(
        ReadAddress[7]), .QN(n654) );
  DFFR_X2 ReadAddress_reg_5_ ( .D(n759), .CK(clock), .RN(n644), .Q(
        ReadAddress[5]) );
  DFFR_X2 ReadAddress_reg_3_ ( .D(n761), .CK(clock), .RN(reset_n), .Q(
        ReadAddress[3]) );
  DFFR_X2 ReadAddress_reg_1_ ( .D(n763), .CK(clock), .RN(reset_n), .Q(
        ReadAddress[1]) );
  AND3_X4 U123 ( .A1(n744), .A2(U6_DATA1_1), .A3(n630), .ZN(n619) );
  AND3_X4 U124 ( .A1(U6_DATA1_1), .A2(U6_DATA1_3), .A3(n630), .ZN(n620) );
  AND2_X4 U125 ( .A1(n632), .A2(n744), .ZN(n621) );
  AND2_X4 U126 ( .A1(n632), .A2(U6_DATA1_3), .ZN(n622) );
  AND2_X4 U127 ( .A1(n633), .A2(n744), .ZN(n623) );
  AND2_X4 U128 ( .A1(n633), .A2(U6_DATA1_3), .ZN(n624) );
  AND2_X4 U129 ( .A1(n744), .A2(n745), .ZN(n625) );
  AND3_X4 U130 ( .A1(n747), .A2(n744), .A3(n746), .ZN(n626) );
  AND3_X4 U131 ( .A1(n747), .A2(U6_DATA1_3), .A3(n746), .ZN(n627) );
  AND2_X4 U132 ( .A1(n745), .A2(U6_DATA1_3), .ZN(n628) );
  AND2_X2 U133 ( .A1(n742), .A2(n741), .ZN(n630) );
  AND3_X4 U134 ( .A1(U6_DATA1_0), .A2(n741), .A3(U6_DATA1_1), .ZN(n631) );
  AND3_X4 U135 ( .A1(n742), .A2(n739), .A3(n746), .ZN(n632) );
  AND2_X4 U136 ( .A1(n747), .A2(n741), .ZN(n633) );
  NOR4_X2 U137 ( .A1(ReadAddress[10]), .A2(ReadAddress[8]), .A3(
        ReadAddress[13]), .A4(n727), .ZN(n656) );
  OAI22_X1 U138 ( .A1(n666), .A2(n725), .B1(n665), .B2(n629), .ZN(n762) );
  NAND3_X2 U139 ( .A1(ReadAddress[4]), .A2(ReadAddress[3]), .A3(n670), .ZN(
        n676) );
  NAND3_X2 U140 ( .A1(ReadAddress[10]), .A2(ReadAddress[9]), .A3(n699), .ZN(
        n702) );
  NAND3_X2 U141 ( .A1(ReadAddress[6]), .A2(ReadAddress[5]), .A3(n679), .ZN(
        n712) );
  MUX2_X1 U142 ( .A(n682), .B(n680), .S(ReadAddress[5]), .Z(n684) );
  NAND3_X1 U144 ( .A1(ReadAddress[1]), .A2(ReadAddress[0]), .A3(ReadAddress[2]), .ZN(n667) );
  OAI22_X1 U145 ( .A1(n725), .A2(n717), .B1(n716), .B2(n727), .ZN(n750) );
  AND2_X4 U146 ( .A1(ReadAddress[12]), .A2(ReadAddress[11]), .ZN(n640) );
  NAND4_X2 U147 ( .A1(ReadAddress[7]), .A2(ReadAddress[9]), .A3(n640), .A4(
        n715), .ZN(n732) );
  MUX2_X1 U149 ( .A(n713), .B(n695), .S(ReadAddress[9]), .Z(n698) );
  MUX2_X1 U150 ( .A(n714), .B(n687), .S(ReadAddress[7]), .Z(n690) );
  NAND3_X1 U151 ( .A1(ReadAddress[8]), .A2(ReadAddress[7]), .A3(n691), .ZN(
        n694) );
  INV_X4 U154 ( .A(n650), .ZN(n645) );
  INV_X4 U155 ( .A(n650), .ZN(n649) );
  INV_X4 U156 ( .A(n650), .ZN(n648) );
  INV_X4 U157 ( .A(n650), .ZN(n647) );
  INV_X4 U159 ( .A(n650), .ZN(n646) );
  INV_X4 U160 ( .A(n650), .ZN(n644) );
  INV_X4 U161 ( .A(n651), .ZN(n749) );
  AND2_X1 U164 ( .A1(n631), .A2(n744), .ZN(n634) );
  AOI21_X2 U165 ( .B1(n722), .B2(n739), .A(n721), .ZN(n723) );
  AND2_X1 U166 ( .A1(U6_DATA1_1), .A2(n746), .ZN(n635) );
  INV_X4 U167 ( .A(reset_n), .ZN(n650) );
  AOI22_X2 U169 ( .A1(U5_DATA2_0), .A2(n749), .B1(U5_DATA1_0), .B2(n621), .ZN(
        n261) );
  AOI22_X2 U170 ( .A1(U5_DATA10_0), .A2(n634), .B1(U5_DATA9_0), .B2(n622), 
        .ZN(n268) );
  AOI22_X2 U171 ( .A1(U5_DATA2_1), .A2(n749), .B1(U5_DATA1_1), .B2(n621), .ZN(
        n251) );
  AOI22_X2 U172 ( .A1(U5_DATA10_1), .A2(n634), .B1(U5_DATA9_1), .B2(n622), 
        .ZN(n255) );
  AOI22_X2 U174 ( .A1(U5_DATA2_2), .A2(n749), .B1(U5_DATA1_2), .B2(n621), .ZN(
        n241) );
  AOI22_X2 U175 ( .A1(U5_DATA10_2), .A2(n634), .B1(U5_DATA9_2), .B2(n622), 
        .ZN(n245) );
  AOI22_X2 U176 ( .A1(U5_DATA2_3), .A2(n749), .B1(U5_DATA1_3), .B2(n621), .ZN(
        n231) );
  AOI22_X2 U177 ( .A1(U5_DATA10_3), .A2(n634), .B1(U5_DATA9_3), .B2(n622), 
        .ZN(n235) );
  AOI22_X2 U179 ( .A1(U5_DATA2_4), .A2(n749), .B1(U5_DATA1_4), .B2(n621), .ZN(
        n221) );
  AOI22_X2 U180 ( .A1(U5_DATA10_4), .A2(n634), .B1(U5_DATA9_4), .B2(n622), 
        .ZN(n225) );
  AOI22_X2 U181 ( .A1(U5_DATA2_5), .A2(n749), .B1(U5_DATA1_5), .B2(n621), .ZN(
        n211) );
  AOI22_X2 U182 ( .A1(U5_DATA10_5), .A2(n634), .B1(U5_DATA9_5), .B2(n622), 
        .ZN(n215) );
  AOI22_X2 U184 ( .A1(U5_DATA2_6), .A2(n749), .B1(U5_DATA1_6), .B2(n621), .ZN(
        n201) );
  AOI22_X2 U185 ( .A1(U5_DATA10_6), .A2(n634), .B1(U5_DATA9_6), .B2(n622), 
        .ZN(n205) );
  AOI22_X2 U186 ( .A1(U5_DATA2_7), .A2(n749), .B1(U5_DATA1_7), .B2(n621), .ZN(
        n175) );
  AOI22_X2 U187 ( .A1(U5_DATA10_7), .A2(n634), .B1(U5_DATA9_7), .B2(n622), 
        .ZN(n187) );
  AOI22_X2 U189 ( .A1(U5_DATA4_0), .A2(n624), .B1(U5_DATA3_0), .B2(n620), .ZN(
        n262) );
  AOI22_X2 U190 ( .A1(U5_DATA12_0), .A2(n623), .B1(U5_DATA11_0), .B2(n619), 
        .ZN(n269) );
  AOI22_X2 U191 ( .A1(U5_DATA4_1), .A2(n624), .B1(U5_DATA3_1), .B2(n620), .ZN(
        n252) );
  AOI22_X2 U192 ( .A1(U5_DATA12_1), .A2(n623), .B1(U5_DATA11_1), .B2(n619), 
        .ZN(n256) );
  AOI22_X2 U194 ( .A1(U5_DATA4_2), .A2(n624), .B1(U5_DATA3_2), .B2(n620), .ZN(
        n242) );
  AOI22_X2 U195 ( .A1(U5_DATA12_2), .A2(n623), .B1(U5_DATA11_2), .B2(n619), 
        .ZN(n246) );
  AOI22_X2 U196 ( .A1(U5_DATA4_3), .A2(n624), .B1(U5_DATA3_3), .B2(n620), .ZN(
        n232) );
  AOI22_X2 U197 ( .A1(U5_DATA12_3), .A2(n623), .B1(U5_DATA11_3), .B2(n619), 
        .ZN(n236) );
  AOI22_X2 U199 ( .A1(U5_DATA4_4), .A2(n624), .B1(U5_DATA3_4), .B2(n620), .ZN(
        n222) );
  AOI22_X2 U200 ( .A1(U5_DATA12_4), .A2(n623), .B1(U5_DATA11_4), .B2(n619), 
        .ZN(n226) );
  AOI22_X2 U201 ( .A1(U5_DATA4_5), .A2(n624), .B1(U5_DATA3_5), .B2(n620), .ZN(
        n212) );
  AOI22_X2 U202 ( .A1(U5_DATA12_5), .A2(n623), .B1(U5_DATA11_5), .B2(n619), 
        .ZN(n216) );
  AOI22_X2 U204 ( .A1(U5_DATA4_6), .A2(n624), .B1(U5_DATA3_6), .B2(n620), .ZN(
        n202) );
  AOI22_X2 U205 ( .A1(U5_DATA12_6), .A2(n623), .B1(U5_DATA11_6), .B2(n619), 
        .ZN(n206) );
  AOI22_X2 U206 ( .A1(U5_DATA4_7), .A2(n624), .B1(U5_DATA3_7), .B2(n620), .ZN(
        n176) );
  AOI22_X2 U207 ( .A1(U5_DATA12_7), .A2(n623), .B1(U5_DATA11_7), .B2(n619), 
        .ZN(n188) );
  AOI22_X2 U209 ( .A1(U5_DATA8_0), .A2(n627), .B1(U5_DATA7_0), .B2(n636), .ZN(
        n264) );
  AOI22_X2 U210 ( .A1(U5_DATA6_0), .A2(n628), .B1(U5_DATA5_0), .B2(n637), .ZN(
        n263) );
  AOI22_X2 U211 ( .A1(U5_DATA16_0), .A2(n626), .B1(U5_DATA15_0), .B2(n638), 
        .ZN(n271) );
  AOI22_X2 U212 ( .A1(U5_DATA14_0), .A2(n625), .B1(U5_DATA13_0), .B2(n639), 
        .ZN(n270) );
  AOI22_X2 U214 ( .A1(U5_DATA8_1), .A2(n627), .B1(U5_DATA7_1), .B2(n636), .ZN(
        n254) );
  AOI22_X2 U215 ( .A1(U5_DATA6_1), .A2(n628), .B1(U5_DATA5_1), .B2(n637), .ZN(
        n253) );
  AOI22_X2 U216 ( .A1(U5_DATA16_1), .A2(n626), .B1(U5_DATA15_1), .B2(n638), 
        .ZN(n258) );
  AOI22_X2 U217 ( .A1(U5_DATA14_1), .A2(n625), .B1(U5_DATA13_1), .B2(n639), 
        .ZN(n257) );
  AOI22_X2 U218 ( .A1(U5_DATA8_2), .A2(n627), .B1(U5_DATA7_2), .B2(n636), .ZN(
        n244) );
  AOI22_X2 U219 ( .A1(U5_DATA6_2), .A2(n628), .B1(U5_DATA5_2), .B2(n637), .ZN(
        n243) );
  AOI22_X2 U220 ( .A1(U5_DATA16_2), .A2(n626), .B1(U5_DATA15_2), .B2(n638), 
        .ZN(n248) );
  AOI22_X2 U221 ( .A1(U5_DATA14_2), .A2(n625), .B1(U5_DATA13_2), .B2(n639), 
        .ZN(n247) );
  AOI22_X2 U222 ( .A1(U5_DATA8_3), .A2(n627), .B1(U5_DATA7_3), .B2(n636), .ZN(
        n234) );
  AOI22_X2 U223 ( .A1(U5_DATA6_3), .A2(n628), .B1(U5_DATA5_3), .B2(n637), .ZN(
        n233) );
  AOI22_X2 U224 ( .A1(U5_DATA16_3), .A2(n626), .B1(U5_DATA15_3), .B2(n638), 
        .ZN(n238) );
  AOI22_X2 U226 ( .A1(U5_DATA14_3), .A2(n625), .B1(U5_DATA13_3), .B2(n639), 
        .ZN(n237) );
  AOI22_X2 U227 ( .A1(U5_DATA8_4), .A2(n627), .B1(U5_DATA7_4), .B2(n636), .ZN(
        n224) );
  AOI22_X2 U228 ( .A1(U5_DATA6_4), .A2(n628), .B1(U5_DATA5_4), .B2(n637), .ZN(
        n223) );
  AOI22_X2 U229 ( .A1(U5_DATA16_4), .A2(n626), .B1(U5_DATA15_4), .B2(n638), 
        .ZN(n228) );
  AOI22_X2 U230 ( .A1(U5_DATA14_4), .A2(n625), .B1(U5_DATA13_4), .B2(n639), 
        .ZN(n227) );
  AOI22_X2 U231 ( .A1(U5_DATA8_5), .A2(n627), .B1(U5_DATA7_5), .B2(n636), .ZN(
        n214) );
  AOI22_X2 U232 ( .A1(U5_DATA6_5), .A2(n628), .B1(U5_DATA5_5), .B2(n637), .ZN(
        n213) );
  AOI22_X2 U233 ( .A1(U5_DATA16_5), .A2(n626), .B1(U5_DATA15_5), .B2(n638), 
        .ZN(n218) );
  AOI22_X2 U234 ( .A1(U5_DATA14_5), .A2(n625), .B1(U5_DATA13_5), .B2(n639), 
        .ZN(n217) );
  AOI22_X2 U235 ( .A1(U5_DATA8_6), .A2(n627), .B1(U5_DATA7_6), .B2(n636), .ZN(
        n204) );
  AOI22_X2 U236 ( .A1(U5_DATA6_6), .A2(n628), .B1(U5_DATA5_6), .B2(n637), .ZN(
        n203) );
  AOI22_X2 U237 ( .A1(U5_DATA16_6), .A2(n626), .B1(U5_DATA15_6), .B2(n638), 
        .ZN(n208) );
  AOI22_X2 U238 ( .A1(U5_DATA14_6), .A2(n625), .B1(U5_DATA13_6), .B2(n639), 
        .ZN(n207) );
  AOI22_X2 U239 ( .A1(U5_DATA8_7), .A2(n627), .B1(U5_DATA7_7), .B2(n636), .ZN(
        n178) );
  AOI22_X2 U240 ( .A1(U5_DATA6_7), .A2(n628), .B1(U5_DATA5_7), .B2(n637), .ZN(
        n177) );
  AOI22_X2 U241 ( .A1(U5_DATA16_7), .A2(n626), .B1(U5_DATA15_7), .B2(n638), 
        .ZN(n190) );
  AOI22_X2 U242 ( .A1(U5_DATA14_7), .A2(n625), .B1(U5_DATA13_7), .B2(n639), 
        .ZN(n189) );
  AND3_X2 U243 ( .A1(U6_DATA1_3), .A2(n742), .A3(n635), .ZN(n636) );
  AND3_X2 U244 ( .A1(n739), .A2(U6_DATA1_3), .A3(n630), .ZN(n637) );
  AND3_X2 U245 ( .A1(n744), .A2(n742), .A3(n635), .ZN(n638) );
  AND3_X2 U246 ( .A1(n744), .A2(n739), .A3(n630), .ZN(n639) );
  OAI21_X1 U247 ( .B1(n660), .B2(n716), .A(n661), .ZN(n281) );
  INV_X4 U248 ( .A(start), .ZN(n643) );
  NAND2_X4 U249 ( .A1(n659), .A2(n658), .ZN(n725) );
  NAND2_X2 U250 ( .A1(n631), .A2(U6_DATA1_3), .ZN(n651) );
  NAND2_X2 U251 ( .A1(start), .A2(n651), .ZN(n726) );
  NAND2_X2 U252 ( .A1(start), .A2(n749), .ZN(n728) );
  INV_X4 U253 ( .A(n728), .ZN(n659) );
  NOR4_X2 U254 ( .A1(n654), .A2(n653), .A3(ReadAddress[12]), .A4(n652), .ZN(
        n655) );
  INV_X4 U255 ( .A(n667), .ZN(n670) );
  INV_X4 U256 ( .A(n676), .ZN(n679) );
  INV_X4 U257 ( .A(n712), .ZN(n691) );
  NAND3_X2 U258 ( .A1(n656), .A2(n655), .A3(n691), .ZN(n658) );
  INV_X4 U259 ( .A(n658), .ZN(n657) );
  NAND2_X2 U260 ( .A1(n659), .A2(n657), .ZN(n748) );
  NAND2_X2 U261 ( .A1(n726), .A2(n748), .ZN(n730) );
  INV_X4 U262 ( .A(n730), .ZN(n716) );
  INV_X4 U263 ( .A(n725), .ZN(n734) );
  NAND2_X2 U264 ( .A1(n734), .A2(n660), .ZN(n661) );
  NOR2_X2 U265 ( .A1(n660), .A2(n725), .ZN(n662) );
  NAND2_X2 U266 ( .A1(n716), .A2(n661), .ZN(n664) );
  MUX2_X2 U267 ( .A(n662), .B(n664), .S(ReadAddress[1]), .Z(n763) );
  NAND2_X2 U268 ( .A1(ReadAddress[0]), .A2(n629), .ZN(n663) );
  MUX2_X2 U269 ( .A(n629), .B(n663), .S(ReadAddress[1]), .Z(n666) );
  INV_X4 U270 ( .A(n664), .ZN(n665) );
  NOR2_X2 U271 ( .A1(n667), .A2(n725), .ZN(n669) );
  NAND2_X2 U272 ( .A1(n734), .A2(n667), .ZN(n668) );
  NAND2_X2 U273 ( .A1(n716), .A2(n668), .ZN(n672) );
  MUX2_X2 U274 ( .A(n669), .B(n672), .S(ReadAddress[3]), .Z(n761) );
  NAND2_X2 U275 ( .A1(n670), .A2(n673), .ZN(n671) );
  MUX2_X2 U276 ( .A(n673), .B(n671), .S(ReadAddress[3]), .Z(n675) );
  INV_X4 U277 ( .A(n672), .ZN(n674) );
  OAI22_X2 U278 ( .A1(n675), .A2(n725), .B1(n674), .B2(n673), .ZN(n760) );
  NOR2_X2 U279 ( .A1(n676), .A2(n725), .ZN(n678) );
  NAND2_X2 U280 ( .A1(n734), .A2(n676), .ZN(n677) );
  NAND2_X2 U281 ( .A1(n716), .A2(n677), .ZN(n681) );
  MUX2_X2 U282 ( .A(n678), .B(n681), .S(ReadAddress[5]), .Z(n759) );
  NAND2_X2 U283 ( .A1(n679), .A2(n682), .ZN(n680) );
  INV_X4 U292 ( .A(n681), .ZN(n683) );
  OAI22_X2 U293 ( .A1(n684), .A2(n725), .B1(n683), .B2(n682), .ZN(n758) );
  NOR2_X2 U294 ( .A1(n712), .A2(n725), .ZN(n686) );
  NAND2_X2 U295 ( .A1(n734), .A2(n712), .ZN(n685) );
  NAND2_X2 U296 ( .A1(n716), .A2(n685), .ZN(n688) );
  MUX2_X2 U297 ( .A(n686), .B(n688), .S(ReadAddress[7]), .Z(n757) );
  NAND2_X2 U298 ( .A1(n691), .A2(n714), .ZN(n687) );
  INV_X4 U299 ( .A(n688), .ZN(n689) );
  OAI22_X2 U300 ( .A1(n690), .A2(n725), .B1(n689), .B2(n714), .ZN(n756) );
  NOR2_X2 U301 ( .A1(n725), .A2(n694), .ZN(n693) );
  NAND2_X2 U302 ( .A1(n734), .A2(n694), .ZN(n692) );
  NAND2_X2 U303 ( .A1(n716), .A2(n692), .ZN(n696) );
  MUX2_X2 U304 ( .A(n693), .B(n696), .S(ReadAddress[9]), .Z(n755) );
  INV_X4 U305 ( .A(n694), .ZN(n699) );
  NAND2_X2 U306 ( .A1(n699), .A2(n713), .ZN(n695) );
  INV_X4 U307 ( .A(n696), .ZN(n697) );
  OAI22_X2 U308 ( .A1(n698), .A2(n725), .B1(n697), .B2(n713), .ZN(n754) );
  NOR2_X2 U309 ( .A1(n725), .A2(n702), .ZN(n701) );
  NAND2_X2 U310 ( .A1(n734), .A2(n702), .ZN(n700) );
  NAND2_X2 U311 ( .A1(n716), .A2(n700), .ZN(n704) );
  MUX2_X2 U312 ( .A(n701), .B(n704), .S(ReadAddress[11]), .Z(n753) );
  INV_X4 U313 ( .A(n702), .ZN(n708) );
  NAND2_X2 U314 ( .A1(n708), .A2(n705), .ZN(n703) );
  MUX2_X2 U315 ( .A(n705), .B(n703), .S(ReadAddress[11]), .Z(n707) );
  INV_X4 U316 ( .A(n704), .ZN(n706) );
  OAI22_X2 U317 ( .A1(n707), .A2(n725), .B1(n706), .B2(n705), .ZN(n752) );
  NAND2_X2 U318 ( .A1(n708), .A2(n640), .ZN(n709) );
  XOR2_X2 U319 ( .A(n709), .B(ReadAddress[13]), .Z(n710) );
  OAI22_X2 U320 ( .A1(n725), .A2(n710), .B1(n716), .B2(n711), .ZN(n751) );
  NOR4_X2 U321 ( .A1(n714), .A2(n713), .A3(n712), .A4(n711), .ZN(n715) );
  XOR2_X2 U322 ( .A(n732), .B(ReadAddress[14]), .Z(n717) );
  INV_X4 U323 ( .A(n726), .ZN(n722) );
  NAND2_X2 U324 ( .A1(n722), .A2(n742), .ZN(n718) );
  NAND2_X2 U325 ( .A1(n748), .A2(n718), .ZN(U3_U5_Z_0) );
  NAND2_X2 U326 ( .A1(n722), .A2(n742), .ZN(n719) );
  NAND2_X2 U327 ( .A1(n719), .A2(n748), .ZN(n721) );
  INV_X4 U328 ( .A(n721), .ZN(n720) );
  NAND2_X2 U329 ( .A1(n739), .A2(U6_DATA1_0), .ZN(n740) );
  OAI22_X2 U330 ( .A1(n739), .A2(n720), .B1(n740), .B2(n726), .ZN(U3_U5_Z_1)
         );
  NAND2_X2 U331 ( .A1(U6_DATA1_0), .A2(n635), .ZN(n743) );
  OAI22_X2 U332 ( .A1(n743), .A2(n726), .B1(n746), .B2(n723), .ZN(U3_U5_Z_2)
         );
  NOR2_X2 U333 ( .A1(U6_DATA1_3), .A2(n631), .ZN(n724) );
  OAI22_X2 U334 ( .A1(n724), .A2(n726), .B1(n723), .B2(n744), .ZN(U3_U5_Z_3)
         );
  NAND2_X2 U335 ( .A1(n726), .A2(n725), .ZN(U3_U3_Z_0) );
  NAND3_X2 U336 ( .A1(output_base_offset), .A2(n728), .A3(n726), .ZN(n738) );
  NOR2_X2 U337 ( .A1(n727), .A2(n732), .ZN(n729) );
  NOR2_X2 U338 ( .A1(n729), .A2(n728), .ZN(n731) );
  NOR2_X2 U339 ( .A1(n731), .A2(n730), .ZN(n736) );
  INV_X4 U340 ( .A(n732), .ZN(n733) );
  NAND3_X2 U341 ( .A1(n734), .A2(ReadAddress[14]), .A3(n733), .ZN(n735) );
  MUX2_X2 U342 ( .A(n736), .B(n735), .S(n147), .Z(n737) );
  NAND2_X2 U343 ( .A1(n738), .A2(n737), .ZN(n280) );
  INV_X4 U344 ( .A(n740), .ZN(n747) );
  INV_X4 U345 ( .A(n743), .ZN(n745) );
  INV_X4 U346 ( .A(n748), .ZN(U3_U4_Z_0) );
  INV_X8 U152 ( .A(n643), .ZN(n641) );
  INV_X8 U162 ( .A(n643), .ZN(n642) );
endmodule


module Output_Fetch_Cdf ( clock, reset_n, ReadBus, ReadAddress, DataIn, 
        DataOut, StartIn, StartOut, output_base_offset );
  input [127:0] ReadBus;
  output [15:0] ReadAddress;
  input [7:0] DataIn;
  output [19:0] DataOut;
  input clock, reset_n, StartIn, output_base_offset;
  output StartOut;

  assign ReadAddress[14] = 1'b0;
  assign ReadAddress[13] = 1'b0;
  assign ReadAddress[12] = 1'b0;
  assign ReadAddress[11] = 1'b0;
  assign ReadAddress[10] = 1'b0;
  assign ReadAddress[9] = 1'b0;
  assign ReadAddress[8] = 1'b0;

  DFF_X1 DataOut_reg_19_ ( .D(ReadBus[19]), .CK(clock), .Q(DataOut[19]) );
  DFF_X1 DataOut_reg_18_ ( .D(ReadBus[18]), .CK(clock), .Q(DataOut[18]) );
  DFF_X1 DataOut_reg_17_ ( .D(ReadBus[17]), .CK(clock), .Q(DataOut[17]) );
  DFF_X1 DataOut_reg_16_ ( .D(ReadBus[16]), .CK(clock), .Q(DataOut[16]) );
  DFF_X1 DataOut_reg_15_ ( .D(ReadBus[15]), .CK(clock), .Q(DataOut[15]) );
  DFF_X1 DataOut_reg_14_ ( .D(ReadBus[14]), .CK(clock), .Q(DataOut[14]) );
  DFF_X1 DataOut_reg_13_ ( .D(ReadBus[13]), .CK(clock), .Q(DataOut[13]) );
  DFF_X1 DataOut_reg_12_ ( .D(ReadBus[12]), .CK(clock), .Q(DataOut[12]) );
  DFF_X1 DataOut_reg_11_ ( .D(ReadBus[11]), .CK(clock), .Q(DataOut[11]) );
  DFF_X1 DataOut_reg_10_ ( .D(ReadBus[10]), .CK(clock), .Q(DataOut[10]) );
  DFF_X1 DataOut_reg_8_ ( .D(ReadBus[8]), .CK(clock), .Q(DataOut[8]) );
  DFF_X1 DataOut_reg_7_ ( .D(ReadBus[7]), .CK(clock), .Q(DataOut[7]) );
  DFF_X1 DataOut_reg_6_ ( .D(ReadBus[6]), .CK(clock), .Q(DataOut[6]) );
  DFF_X1 DataOut_reg_5_ ( .D(ReadBus[5]), .CK(clock), .Q(DataOut[5]) );
  DFF_X1 DataOut_reg_4_ ( .D(ReadBus[4]), .CK(clock), .Q(DataOut[4]) );
  DFF_X1 DataOut_reg_3_ ( .D(ReadBus[3]), .CK(clock), .Q(DataOut[3]) );
  DFF_X1 DataOut_reg_2_ ( .D(ReadBus[2]), .CK(clock), .Q(DataOut[2]) );
  DFF_X1 DataOut_reg_1_ ( .D(ReadBus[1]), .CK(clock), .Q(DataOut[1]) );
  DFF_X1 DataOut_reg_0_ ( .D(ReadBus[0]), .CK(clock), .Q(DataOut[0]) );
  DFF_X2 DataOut_reg_9_ ( .D(ReadBus[9]), .CK(clock), .Q(DataOut[9]) );
  DFFR_X2 StartOut_reg ( .D(StartIn), .CK(clock), .RN(reset_n), .Q(StartOut)
         );
  BUF_X4 U17 ( .A(output_base_offset), .Z(ReadAddress[15]) );
  BUF_X4 U18 ( .A(DataIn[7]), .Z(ReadAddress[7]) );
  BUF_X4 U19 ( .A(DataIn[6]), .Z(ReadAddress[6]) );
  BUF_X4 U20 ( .A(DataIn[5]), .Z(ReadAddress[5]) );
  BUF_X4 U21 ( .A(DataIn[4]), .Z(ReadAddress[4]) );
  BUF_X4 U22 ( .A(DataIn[3]), .Z(ReadAddress[3]) );
  BUF_X4 U23 ( .A(DataIn[2]), .Z(ReadAddress[2]) );
  BUF_X4 U24 ( .A(DataIn[1]), .Z(ReadAddress[1]) );
  BUF_X4 U25 ( .A(DataIn[0]), .Z(ReadAddress[0]) );
endmodule


module Output_TopExpression ( clock, reset_n, DataIn, CdfMin, StartIn, 
        StartOut, DataOut );
  input [19:0] DataIn;
  input [19:0] CdfMin;
  output [27:0] DataOut;
  input clock, reset_n, StartIn;
  output StartOut;
  wire   U4_Z_0, U4_Z_1, U4_Z_2, U4_Z_3, U4_Z_4, U4_Z_5, U4_Z_6, U4_Z_7,
         U4_Z_8, U4_Z_9, U4_Z_10, U4_Z_11, U4_Z_12, U4_Z_13, U4_Z_14, U4_Z_15,
         U4_Z_16, U4_Z_17, U4_Z_18, U4_Z_19, U4_Z_21, U4_Z_22, U4_Z_24,
         U4_Z_26, U4_Z_27, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818;

  DFFR_X1 DataOut_reg_13_ ( .D(U4_Z_13), .CK(clock), .RN(n365), .Q(DataOut[13]) );
  DFFR_X1 DataOut_reg_12_ ( .D(U4_Z_12), .CK(clock), .RN(n365), .Q(DataOut[12]) );
  DFFR_X1 DataOut_reg_11_ ( .D(U4_Z_11), .CK(clock), .RN(n364), .Q(DataOut[11]) );
  DFFR_X1 DataOut_reg_10_ ( .D(U4_Z_10), .CK(clock), .RN(n364), .Q(DataOut[10]) );
  DFFR_X1 DataOut_reg_9_ ( .D(U4_Z_9), .CK(clock), .RN(n364), .Q(DataOut[9])
         );
  DFFR_X1 DataOut_reg_8_ ( .D(U4_Z_8), .CK(clock), .RN(n364), .Q(DataOut[8])
         );
  DFFR_X1 DataOut_reg_7_ ( .D(U4_Z_7), .CK(clock), .RN(n364), .Q(DataOut[7])
         );
  DFFR_X2 DataOut_reg_15_ ( .D(U4_Z_15), .CK(clock), .RN(reset_n), .Q(
        DataOut[15]) );
  DFFR_X2 DataOut_reg_17_ ( .D(U4_Z_17), .CK(clock), .RN(n365), .Q(DataOut[17]) );
  DFFR_X2 DataOut_reg_19_ ( .D(U4_Z_19), .CK(clock), .RN(n365), .Q(DataOut[19]) );
  DFFR_X2 DataOut_reg_18_ ( .D(U4_Z_18), .CK(clock), .RN(n365), .Q(DataOut[18]) );
  DFFR_X2 DataOut_reg_24_ ( .D(U4_Z_24), .CK(clock), .RN(n365), .Q(DataOut[24]) );
  DFFR_X2 DataOut_reg_22_ ( .D(U4_Z_22), .CK(clock), .RN(n365), .Q(DataOut[22]) );
  DFFR_X2 DataOut_reg_23_ ( .D(n817), .CK(clock), .RN(n365), .Q(DataOut[23])
         );
  DFFR_X2 DataOut_reg_21_ ( .D(U4_Z_21), .CK(clock), .RN(n365), .Q(DataOut[21]) );
  DFFR_X2 DataOut_reg_16_ ( .D(U4_Z_16), .CK(clock), .RN(n365), .Q(DataOut[16]) );
  DFFR_X1 DataOut_reg_27_ ( .D(U4_Z_27), .CK(clock), .RN(n364), .Q(DataOut[27]) );
  DFFR_X1 DataOut_reg_26_ ( .D(U4_Z_26), .CK(clock), .RN(n365), .Q(DataOut[26]) );
  DFFR_X1 DataOut_reg_25_ ( .D(n818), .CK(clock), .RN(n365), .Q(DataOut[25])
         );
  DFFR_X2 StartOut_reg ( .D(StartIn), .CK(clock), .RN(n364), .Q(StartOut) );
  DFFR_X2 DataOut_reg_0_ ( .D(U4_Z_0), .CK(clock), .RN(n364), .Q(DataOut[0])
         );
  DFFR_X2 DataOut_reg_1_ ( .D(U4_Z_1), .CK(clock), .RN(n364), .Q(DataOut[1])
         );
  DFFR_X2 DataOut_reg_5_ ( .D(U4_Z_5), .CK(clock), .RN(n364), .Q(DataOut[5])
         );
  DFFR_X2 DataOut_reg_2_ ( .D(U4_Z_2), .CK(clock), .RN(n364), .Q(DataOut[2])
         );
  DFFR_X2 DataOut_reg_4_ ( .D(U4_Z_4), .CK(clock), .RN(n364), .Q(DataOut[4])
         );
  DFFR_X2 DataOut_reg_6_ ( .D(U4_Z_6), .CK(clock), .RN(n364), .Q(DataOut[6])
         );
  DFFR_X2 DataOut_reg_3_ ( .D(U4_Z_3), .CK(clock), .RN(reset_n), .Q(DataOut[3]) );
  DFFR_X2 DataOut_reg_14_ ( .D(U4_Z_14), .CK(clock), .RN(reset_n), .Q(
        DataOut[14]) );
  DFFR_X1 DataOut_reg_20_ ( .D(n816), .CK(clock), .RN(n365), .Q(DataOut[20])
         );
  INV_X4 U3 ( .A(n399), .ZN(n242) );
  INV_X1 U4 ( .A(n425), .ZN(n428) );
  INV_X1 U5 ( .A(n810), .ZN(n159) );
  INV_X2 U6 ( .A(n758), .ZN(n160) );
  NAND2_X1 U7 ( .A1(n731), .A2(n780), .ZN(n741) );
  INV_X2 U8 ( .A(n660), .ZN(n161) );
  INV_X2 U9 ( .A(n673), .ZN(n660) );
  NAND2_X1 U10 ( .A1(n186), .A2(n810), .ZN(n778) );
  OAI221_X2 U11 ( .B1(n753), .B2(n768), .C1(n806), .C2(n748), .A(StartIn), 
        .ZN(n749) );
  NAND2_X4 U12 ( .A1(n666), .A2(n681), .ZN(n720) );
  NOR2_X1 U13 ( .A1(n724), .A2(n719), .ZN(n699) );
  INV_X2 U14 ( .A(n389), .ZN(n162) );
  INV_X4 U15 ( .A(n162), .ZN(n163) );
  INV_X4 U16 ( .A(n807), .ZN(n806) );
  INV_X4 U17 ( .A(n620), .ZN(n241) );
  NAND3_X2 U18 ( .A1(n743), .A2(n814), .A3(n742), .ZN(n208) );
  NAND2_X2 U19 ( .A1(n549), .A2(n548), .ZN(n164) );
  NAND2_X2 U20 ( .A1(n296), .A2(n297), .ZN(n165) );
  NAND2_X2 U21 ( .A1(n633), .A2(n608), .ZN(n168) );
  NAND2_X2 U22 ( .A1(n166), .A2(n167), .ZN(n169) );
  NAND2_X2 U23 ( .A1(n168), .A2(n169), .ZN(n263) );
  INV_X2 U24 ( .A(n633), .ZN(n166) );
  INV_X4 U25 ( .A(n608), .ZN(n167) );
  INV_X1 U26 ( .A(n607), .ZN(n608) );
  OR2_X2 U27 ( .A1(n263), .A2(n610), .ZN(n297) );
  INV_X4 U28 ( .A(n263), .ZN(n622) );
  NAND2_X2 U29 ( .A1(n678), .A2(n345), .ZN(n606) );
  INV_X4 U30 ( .A(n564), .ZN(n286) );
  AND2_X2 U31 ( .A1(n543), .A2(n342), .ZN(n170) );
  INV_X2 U32 ( .A(DataIn[3]), .ZN(n384) );
  INV_X4 U33 ( .A(n546), .ZN(n221) );
  AND2_X1 U34 ( .A1(n412), .A2(n454), .ZN(n171) );
  INV_X2 U35 ( .A(n615), .ZN(n624) );
  NAND2_X4 U36 ( .A1(n623), .A2(n215), .ZN(n308) );
  AND2_X4 U37 ( .A1(n759), .A2(n760), .ZN(n172) );
  INV_X1 U38 ( .A(n388), .ZN(n173) );
  INV_X1 U39 ( .A(n173), .ZN(n174) );
  NOR3_X2 U40 ( .A1(n266), .A2(n267), .A3(n315), .ZN(n175) );
  NOR3_X2 U41 ( .A1(n266), .A2(n267), .A3(n315), .ZN(n511) );
  INV_X1 U42 ( .A(n261), .ZN(n552) );
  NAND2_X4 U43 ( .A1(n488), .A2(n280), .ZN(n518) );
  INV_X2 U44 ( .A(n734), .ZN(n659) );
  INV_X1 U45 ( .A(n306), .ZN(n307) );
  AND2_X2 U46 ( .A1(n382), .A2(n174), .ZN(n237) );
  INV_X1 U47 ( .A(n363), .ZN(n176) );
  INV_X2 U48 ( .A(n176), .ZN(n177) );
  NAND2_X4 U49 ( .A1(n305), .A2(n170), .ZN(n599) );
  OR2_X1 U50 ( .A1(n240), .A2(n235), .ZN(n178) );
  OR2_X1 U51 ( .A1(n434), .A2(n433), .ZN(n179) );
  NAND3_X2 U52 ( .A1(n178), .A2(n179), .A3(n432), .ZN(n620) );
  NAND2_X1 U53 ( .A1(n412), .A2(n454), .ZN(n230) );
  NAND2_X2 U54 ( .A1(n514), .A2(n513), .ZN(n515) );
  NAND2_X2 U55 ( .A1(n172), .A2(n758), .ZN(n763) );
  NOR2_X1 U56 ( .A1(n754), .A2(n753), .ZN(n760) );
  NAND2_X1 U57 ( .A1(n770), .A2(n254), .ZN(n761) );
  INV_X2 U58 ( .A(n769), .ZN(n772) );
  INV_X1 U59 ( .A(n412), .ZN(n416) );
  NAND2_X2 U60 ( .A1(n609), .A2(n637), .ZN(n702) );
  INV_X2 U61 ( .A(n307), .ZN(n184) );
  AOI21_X2 U62 ( .B1(n708), .B2(n784), .A(n672), .ZN(n671) );
  AND2_X2 U63 ( .A1(n731), .A2(n711), .ZN(n180) );
  INV_X4 U64 ( .A(n759), .ZN(n256) );
  INV_X4 U65 ( .A(n739), .ZN(n740) );
  AND2_X4 U66 ( .A1(n814), .A2(n180), .ZN(n181) );
  AND2_X1 U67 ( .A1(n707), .A2(n721), .ZN(n182) );
  INV_X4 U68 ( .A(n580), .ZN(n270) );
  INV_X4 U69 ( .A(n788), .ZN(n795) );
  INV_X2 U70 ( .A(n575), .ZN(n356) );
  INV_X2 U71 ( .A(n324), .ZN(n400) );
  INV_X4 U72 ( .A(DataIn[8]), .ZN(n348) );
  INV_X4 U73 ( .A(n426), .ZN(n442) );
  OAI22_X2 U74 ( .A1(n592), .A2(n610), .B1(n759), .B2(n591), .ZN(n604) );
  XNOR2_X2 U75 ( .A(n227), .B(n184), .ZN(n183) );
  INV_X4 U76 ( .A(n183), .ZN(n226) );
  NAND2_X2 U77 ( .A1(n425), .A2(n200), .ZN(n223) );
  NOR2_X2 U78 ( .A1(n778), .A2(n185), .ZN(n278) );
  OR2_X1 U79 ( .A1(n780), .A2(n781), .ZN(n185) );
  NOR3_X2 U80 ( .A1(n277), .A2(n278), .A3(n777), .ZN(U4_Z_24) );
  AND2_X1 U81 ( .A1(n778), .A2(n780), .ZN(n277) );
  NAND2_X2 U82 ( .A1(n233), .A2(n190), .ZN(n734) );
  XNOR2_X2 U83 ( .A(n659), .B(n339), .ZN(n635) );
  INV_X2 U84 ( .A(n677), .ZN(U4_Z_18) );
  NAND2_X1 U85 ( .A1(n781), .A2(n780), .ZN(n776) );
  NAND2_X2 U86 ( .A1(n744), .A2(n208), .ZN(n786) );
  INV_X2 U87 ( .A(n254), .ZN(n783) );
  NAND2_X2 U88 ( .A1(n293), .A2(n810), .ZN(n812) );
  INV_X2 U89 ( .A(n255), .ZN(n658) );
  NAND2_X1 U90 ( .A1(n809), .A2(n815), .ZN(n794) );
  NOR3_X1 U91 ( .A1(n815), .A2(n809), .A3(n814), .ZN(n813) );
  NAND2_X1 U92 ( .A1(n320), .A2(n321), .ZN(n244) );
  INV_X4 U93 ( .A(n417), .ZN(n468) );
  NAND2_X4 U94 ( .A1(n276), .A2(n452), .ZN(n409) );
  NAND2_X2 U95 ( .A1(n488), .A2(n280), .ZN(n252) );
  NAND2_X1 U96 ( .A1(n757), .A2(n795), .ZN(n186) );
  XNOR2_X1 U97 ( .A(n252), .B(n351), .ZN(n187) );
  XNOR2_X2 U98 ( .A(n500), .B(n260), .ZN(n351) );
  NAND2_X2 U99 ( .A1(n757), .A2(n795), .ZN(n254) );
  CLKBUF_X3 U100 ( .A(n470), .Z(n188) );
  INV_X4 U101 ( .A(n765), .ZN(U4_Z_22) );
  NAND2_X2 U102 ( .A1(n175), .A2(n510), .ZN(n189) );
  NAND2_X2 U103 ( .A1(n511), .A2(n510), .ZN(n544) );
  NAND2_X2 U104 ( .A1(n164), .A2(n766), .ZN(n581) );
  NAND2_X1 U105 ( .A1(n631), .A2(n308), .ZN(n190) );
  AND2_X2 U106 ( .A1(n503), .A2(n205), .ZN(n267) );
  OR2_X1 U107 ( .A1(n300), .A2(n299), .ZN(n654) );
  NOR2_X2 U108 ( .A1(n653), .A2(n360), .ZN(n299) );
  XOR2_X1 U109 ( .A(n226), .B(n476), .Z(n370) );
  NAND2_X1 U110 ( .A1(n226), .A2(StartIn), .ZN(n372) );
  INV_X4 U111 ( .A(n198), .ZN(n582) );
  NAND2_X4 U112 ( .A1(n578), .A2(n579), .ZN(n563) );
  INV_X4 U113 ( .A(n374), .ZN(n306) );
  INV_X2 U114 ( .A(n407), .ZN(n201) );
  INV_X8 U115 ( .A(CdfMin[5]), .ZN(n407) );
  NAND2_X1 U116 ( .A1(n249), .A2(n217), .ZN(n191) );
  NAND2_X2 U117 ( .A1(n379), .A2(n216), .ZN(n192) );
  NAND2_X2 U118 ( .A1(n191), .A2(n192), .ZN(n469) );
  INV_X1 U119 ( .A(n379), .ZN(n249) );
  INV_X1 U120 ( .A(n216), .ZN(n217) );
  INV_X1 U121 ( .A(n471), .ZN(n460) );
  AND2_X4 U122 ( .A1(n258), .A2(n563), .ZN(n331) );
  NAND3_X2 U123 ( .A1(n224), .A2(n193), .A3(n194), .ZN(n281) );
  NAND2_X1 U124 ( .A1(n559), .A2(n558), .ZN(n193) );
  NAND2_X1 U125 ( .A1(n561), .A2(n560), .ZN(n194) );
  NAND2_X1 U126 ( .A1(n440), .A2(DataIn[7]), .ZN(n196) );
  NAND2_X2 U127 ( .A1(n195), .A2(n451), .ZN(n197) );
  NAND2_X2 U128 ( .A1(n196), .A2(n197), .ZN(n350) );
  INV_X2 U129 ( .A(n440), .ZN(n195) );
  OAI22_X2 U130 ( .A1(n545), .A2(n207), .B1(n614), .B2(n548), .ZN(n198) );
  NOR2_X1 U131 ( .A1(n487), .A2(DataIn[9]), .ZN(n199) );
  NOR2_X2 U132 ( .A1(n487), .A2(DataIn[9]), .ZN(n246) );
  INV_X4 U133 ( .A(n442), .ZN(n200) );
  INV_X2 U134 ( .A(n548), .ZN(n550) );
  NAND3_X2 U135 ( .A1(n405), .A2(n548), .A3(n221), .ZN(n435) );
  NAND2_X2 U136 ( .A1(n211), .A2(n200), .ZN(n413) );
  INV_X1 U137 ( .A(n243), .ZN(n202) );
  INV_X2 U138 ( .A(n242), .ZN(n243) );
  NAND2_X2 U139 ( .A1(n581), .A2(n616), .ZN(n203) );
  NAND2_X2 U140 ( .A1(n721), .A2(n562), .ZN(n222) );
  NAND2_X2 U141 ( .A1(n549), .A2(n548), .ZN(n257) );
  NAND2_X1 U142 ( .A1(n310), .A2(n494), .ZN(n204) );
  OR2_X1 U143 ( .A1(n582), .A2(n563), .ZN(n322) );
  NAND2_X1 U144 ( .A1(n624), .A2(n551), .ZN(n577) );
  INV_X1 U145 ( .A(n567), .ZN(n258) );
  XOR2_X1 U146 ( .A(n201), .B(n408), .Z(n396) );
  NAND2_X2 U147 ( .A1(CdfMin[5]), .A2(n408), .ZN(n453) );
  NAND3_X2 U148 ( .A1(n323), .A2(n322), .A3(n273), .ZN(n261) );
  OR2_X1 U149 ( .A1(n582), .A2(n222), .ZN(n323) );
  NOR2_X1 U150 ( .A1(n502), .A2(n199), .ZN(n205) );
  NOR2_X1 U151 ( .A1(n502), .A2(n199), .ZN(n206) );
  INV_X2 U152 ( .A(n213), .ZN(n330) );
  NOR3_X4 U153 ( .A1(n326), .A2(n327), .A3(n328), .ZN(n207) );
  INV_X8 U154 ( .A(n207), .ZN(n766) );
  INV_X1 U155 ( .A(n466), .ZN(n209) );
  INV_X1 U156 ( .A(n209), .ZN(n210) );
  INV_X2 U157 ( .A(n444), .ZN(n211) );
  OR2_X1 U158 ( .A1(n487), .A2(DataIn[9]), .ZN(n212) );
  NAND3_X1 U159 ( .A1(n581), .A2(n222), .A3(n580), .ZN(n213) );
  INV_X1 U160 ( .A(n628), .ZN(n214) );
  INV_X4 U161 ( .A(n214), .ZN(n215) );
  INV_X1 U162 ( .A(n735), .ZN(n233) );
  INV_X1 U163 ( .A(n303), .ZN(n216) );
  INV_X2 U164 ( .A(n533), .ZN(n328) );
  INV_X1 U165 ( .A(n373), .ZN(n218) );
  INV_X4 U166 ( .A(n218), .ZN(n219) );
  NAND2_X2 U167 ( .A1(n368), .A2(n369), .ZN(n373) );
  INV_X4 U168 ( .A(n316), .ZN(n447) );
  INV_X4 U169 ( .A(n614), .ZN(n546) );
  NAND2_X2 U170 ( .A1(n475), .A2(n476), .ZN(n220) );
  NAND2_X2 U171 ( .A1(n241), .A2(n622), .ZN(n628) );
  NAND2_X1 U172 ( .A1(n263), .A2(n620), .ZN(n621) );
  XNOR2_X2 U173 ( .A(n188), .B(n223), .ZN(n548) );
  INV_X2 U174 ( .A(n557), .ZN(n224) );
  OAI211_X4 U175 ( .C1(n261), .C2(n617), .A(n165), .B(n588), .ZN(n618) );
  XOR2_X2 U176 ( .A(n189), .B(n354), .Z(n225) );
  XNOR2_X2 U177 ( .A(DataIn[1]), .B(n369), .ZN(n227) );
  NAND2_X2 U178 ( .A1(n490), .A2(n220), .ZN(n492) );
  NAND2_X2 U179 ( .A1(n565), .A2(n616), .ZN(n568) );
  NAND2_X2 U180 ( .A1(n491), .A2(n226), .ZN(n310) );
  NAND2_X2 U181 ( .A1(n729), .A2(n728), .ZN(n739) );
  NAND2_X2 U182 ( .A1(n641), .A2(n606), .ZN(n609) );
  INV_X1 U183 ( .A(n526), .ZN(n228) );
  INV_X4 U184 ( .A(n228), .ZN(n229) );
  NAND2_X2 U185 ( .A1(n304), .A2(n424), .ZN(n526) );
  INV_X4 U186 ( .A(n264), .ZN(n265) );
  NAND3_X2 U187 ( .A1(n509), .A2(n508), .A3(n507), .ZN(n264) );
  INV_X2 U188 ( .A(n712), .ZN(n714) );
  NAND2_X2 U189 ( .A1(n412), .A2(n454), .ZN(n481) );
  INV_X1 U190 ( .A(n795), .ZN(n231) );
  NAND2_X2 U191 ( .A1(n626), .A2(n238), .ZN(n232) );
  INV_X2 U192 ( .A(n291), .ZN(n657) );
  INV_X1 U193 ( .A(n438), .ZN(n234) );
  INV_X4 U194 ( .A(n234), .ZN(n235) );
  INV_X1 U195 ( .A(n506), .ZN(n236) );
  NAND2_X2 U196 ( .A1(n355), .A2(DataIn[6]), .ZN(n438) );
  AND2_X4 U197 ( .A1(n507), .A2(n245), .ZN(n266) );
  XNOR2_X2 U198 ( .A(n237), .B(n353), .ZN(n614) );
  INV_X2 U199 ( .A(CdfMin[7]), .ZN(n440) );
  INV_X2 U200 ( .A(DataIn[7]), .ZN(n451) );
  BUF_X4 U201 ( .A(n350), .Z(n240) );
  OAI221_X2 U202 ( .B1(n286), .B2(n652), .C1(n232), .C2(n330), .A(n651), .ZN(
        n631) );
  NAND2_X2 U203 ( .A1(n455), .A2(n454), .ZN(n508) );
  NAND2_X1 U204 ( .A1(CdfMin[3]), .A2(n384), .ZN(n386) );
  INV_X2 U205 ( .A(n517), .ZN(n579) );
  INV_X2 U206 ( .A(n381), .ZN(n303) );
  INV_X2 U207 ( .A(n587), .ZN(n238) );
  NAND2_X2 U208 ( .A1(n576), .A2(n616), .ZN(n625) );
  INV_X2 U209 ( .A(n355), .ZN(n304) );
  NAND2_X1 U210 ( .A1(n527), .A2(n526), .ZN(n478) );
  NAND2_X1 U211 ( .A1(n229), .A2(n230), .ZN(n427) );
  NAND2_X1 U212 ( .A1(n217), .A2(n379), .ZN(n239) );
  NAND2_X2 U213 ( .A1(n409), .A2(n453), .ZN(n455) );
  NAND2_X2 U214 ( .A1(DataIn[0]), .A2(n375), .ZN(n368) );
  INV_X4 U215 ( .A(n551), .ZN(n653) );
  OR2_X2 U216 ( .A1(n374), .A2(DataIn[1]), .ZN(n302) );
  NAND2_X2 U217 ( .A1(n490), .A2(n489), .ZN(n512) );
  NAND2_X1 U218 ( .A1(n450), .A2(n449), .ZN(n245) );
  INV_X4 U219 ( .A(CdfMin[9]), .ZN(n487) );
  INV_X2 U220 ( .A(DataIn[9]), .ZN(n484) );
  NAND2_X2 U221 ( .A1(n734), .A2(n181), .ZN(n744) );
  INV_X2 U222 ( .A(n652), .ZN(n359) );
  XNOR2_X1 U223 ( .A(n201), .B(DataIn[5]), .ZN(n402) );
  AND2_X1 U224 ( .A1(n210), .A2(n465), .ZN(n334) );
  NAND2_X2 U225 ( .A1(n208), .A2(n744), .ZN(n247) );
  XNOR2_X2 U226 ( .A(n390), .B(DataIn[3]), .ZN(n353) );
  NOR2_X2 U227 ( .A1(n250), .A2(n251), .ZN(n248) );
  INV_X4 U228 ( .A(n499), .ZN(n502) );
  NAND2_X2 U229 ( .A1(n706), .A2(n182), .ZN(n709) );
  NOR3_X1 U230 ( .A1(n716), .A2(n700), .A3(n699), .ZN(n707) );
  INV_X1 U231 ( .A(n609), .ZN(n602) );
  NAND2_X1 U232 ( .A1(n702), .A2(n701), .ZN(n717) );
  NOR2_X1 U233 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR3_X4 U234 ( .A1(n444), .A2(n443), .A3(n442), .ZN(n448) );
  NOR2_X2 U235 ( .A1(n502), .A2(n501), .ZN(n250) );
  NOR2_X1 U236 ( .A1(CdfMin[10]), .A2(n500), .ZN(n251) );
  XNOR2_X2 U237 ( .A(n306), .B(DataIn[1]), .ZN(n459) );
  NAND2_X2 U238 ( .A1(n356), .A2(n271), .ZN(n320) );
  NAND2_X1 U239 ( .A1(n380), .A2(n239), .ZN(n382) );
  NAND3_X1 U240 ( .A1(n476), .A2(n517), .A3(n183), .ZN(n391) );
  XNOR2_X1 U241 ( .A(n669), .B(n517), .ZN(n495) );
  NOR2_X1 U242 ( .A1(n243), .A2(n400), .ZN(n401) );
  INV_X2 U243 ( .A(n454), .ZN(n443) );
  NAND2_X4 U244 ( .A1(n407), .A2(DataIn[5]), .ZN(n454) );
  NAND2_X1 U245 ( .A1(n367), .A2(CdfMin[0]), .ZN(n301) );
  INV_X2 U246 ( .A(DataIn[0]), .ZN(n367) );
  NAND2_X2 U247 ( .A1(n466), .A2(n465), .ZN(n253) );
  NAND2_X2 U248 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U249 ( .A1(n233), .A2(n656), .ZN(n255) );
  INV_X4 U250 ( .A(n761), .ZN(n758) );
  INV_X1 U251 ( .A(n380), .ZN(n376) );
  INV_X4 U252 ( .A(CdfMin[4]), .ZN(n275) );
  NAND3_X2 U253 ( .A1(n468), .A2(n469), .A3(n470), .ZN(n472) );
  NAND2_X2 U254 ( .A1(n253), .A2(n352), .ZN(n284) );
  NAND2_X1 U255 ( .A1(n175), .A2(n510), .ZN(n298) );
  INV_X4 U256 ( .A(n478), .ZN(n509) );
  NAND2_X2 U257 ( .A1(n504), .A2(n530), .ZN(n477) );
  INV_X2 U258 ( .A(n504), .ZN(n457) );
  NAND2_X2 U259 ( .A1(n530), .A2(n342), .ZN(n313) );
  NAND2_X2 U260 ( .A1(n657), .A2(n656), .ZN(n269) );
  INV_X4 U261 ( .A(n613), .ZN(n567) );
  INV_X1 U262 ( .A(CdfMin[10]), .ZN(n259) );
  INV_X2 U263 ( .A(n259), .ZN(n260) );
  XOR2_X1 U264 ( .A(n305), .B(n347), .Z(n713) );
  OAI22_X1 U265 ( .A1(n331), .A2(n221), .B1(n795), .B2(n653), .ZN(n536) );
  NAND4_X1 U266 ( .A1(n474), .A2(n460), .A3(n614), .A4(n517), .ZN(n462) );
  AND3_X2 U267 ( .A1(n229), .A2(n230), .A3(n527), .ZN(n529) );
  XNOR2_X2 U268 ( .A(n424), .B(n355), .ZN(n415) );
  INV_X1 U269 ( .A(n487), .ZN(n262) );
  INV_X2 U270 ( .A(n271), .ZN(n290) );
  XOR2_X2 U271 ( .A(n276), .B(n452), .Z(n470) );
  NAND2_X2 U272 ( .A1(n389), .A2(n445), .ZN(n288) );
  INV_X1 U273 ( .A(n248), .ZN(n315) );
  NAND2_X2 U274 ( .A1(n459), .A2(n476), .ZN(n471) );
  NAND3_X2 U275 ( .A1(n530), .A2(n509), .A3(n481), .ZN(n294) );
  INV_X1 U276 ( .A(n441), .ZN(n444) );
  NAND4_X4 U277 ( .A1(n697), .A2(n696), .A3(n695), .A4(n694), .ZN(n814) );
  NAND2_X2 U278 ( .A1(n528), .A2(n265), .ZN(n510) );
  INV_X4 U279 ( .A(n497), .ZN(n507) );
  NOR2_X1 U280 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND3_X2 U281 ( .A1(n258), .A2(n580), .A3(n221), .ZN(n551) );
  INV_X1 U282 ( .A(n498), .ZN(n503) );
  NOR2_X2 U283 ( .A1(n566), .A2(n203), .ZN(n570) );
  INV_X1 U284 ( .A(n539), .ZN(n268) );
  INV_X1 U285 ( .A(n281), .ZN(n759) );
  NAND3_X1 U286 ( .A1(n425), .A2(n398), .A3(n394), .ZN(n404) );
  NAND2_X2 U287 ( .A1(n582), .A2(n581), .ZN(n626) );
  INV_X2 U288 ( .A(n467), .ZN(n282) );
  NAND2_X2 U289 ( .A1(n367), .A2(CdfMin[0]), .ZN(n369) );
  INV_X4 U290 ( .A(n678), .ZN(n271) );
  INV_X4 U291 ( .A(n275), .ZN(n276) );
  NAND2_X2 U292 ( .A1(n600), .A2(n599), .ZN(n678) );
  INV_X2 U293 ( .A(n601), .ZN(n645) );
  NOR2_X2 U294 ( .A1(n653), .A2(n615), .ZN(n617) );
  NOR2_X2 U295 ( .A1(n546), .A2(n391), .ZN(n392) );
  NAND2_X2 U296 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X4 U297 ( .A(n770), .ZN(n771) );
  NAND2_X1 U298 ( .A1(n439), .A2(n527), .ZN(n272) );
  NAND2_X2 U299 ( .A1(n439), .A2(n527), .ZN(n450) );
  NAND2_X2 U300 ( .A1(n450), .A2(n449), .ZN(n504) );
  BUF_X4 U301 ( .A(n581), .Z(n273) );
  NOR2_X2 U302 ( .A1(n274), .A2(n783), .ZN(n318) );
  NAND2_X2 U303 ( .A1(n747), .A2(n750), .ZN(n274) );
  XOR2_X1 U304 ( .A(n546), .B(n405), .Z(n383) );
  XNOR2_X2 U305 ( .A(n717), .B(n346), .ZN(n780) );
  INV_X1 U306 ( .A(n501), .ZN(n279) );
  INV_X1 U307 ( .A(n279), .ZN(n280) );
  NOR3_X1 U308 ( .A1(n442), .A2(n415), .A3(n428), .ZN(n414) );
  NAND3_X1 U309 ( .A1(n415), .A2(n413), .A3(n416), .ZN(n420) );
  OAI221_X2 U310 ( .B1(n810), .B2(n746), .C1(n358), .C2(n746), .A(n745), .ZN(
        n816) );
  NAND2_X2 U311 ( .A1(n562), .A2(n721), .ZN(n613) );
  NAND2_X2 U312 ( .A1(n282), .A2(n283), .ZN(n285) );
  NAND2_X2 U313 ( .A1(n284), .A2(n285), .ZN(n490) );
  INV_X1 U314 ( .A(n352), .ZN(n283) );
  XNOR2_X2 U315 ( .A(n348), .B(CdfMin[8]), .ZN(n352) );
  INV_X1 U316 ( .A(n611), .ZN(n571) );
  NOR2_X1 U317 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR3_X1 U318 ( .A1(n226), .A2(n804), .A3(n219), .ZN(n377) );
  NAND2_X1 U319 ( .A1(StartIn), .A2(n219), .ZN(n371) );
  NAND3_X1 U320 ( .A1(n211), .A2(n454), .A3(n414), .ZN(n419) );
  NAND2_X1 U321 ( .A1(n395), .A2(n211), .ZN(n397) );
  NAND2_X2 U322 ( .A1(n445), .A2(n163), .ZN(n287) );
  NAND2_X2 U323 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X2 U324 ( .A1(n325), .A2(n308), .ZN(n362) );
  NAND2_X2 U325 ( .A1(CdfMin[7]), .A2(n451), .ZN(n527) );
  NAND3_X2 U326 ( .A1(n314), .A2(n528), .A3(n529), .ZN(n534) );
  NOR2_X4 U327 ( .A1(n502), .A2(n246), .ZN(n341) );
  INV_X4 U328 ( .A(CdfMin[6]), .ZN(n355) );
  INV_X1 U329 ( .A(n491), .ZN(n289) );
  NAND2_X1 U330 ( .A1(n350), .A2(n235), .ZN(n433) );
  NAND2_X4 U331 ( .A1(n491), .A2(n226), .ZN(n516) );
  INV_X1 U332 ( .A(n626), .ZN(n583) );
  NOR3_X1 U333 ( .A1(n425), .A2(n240), .A3(n427), .ZN(n431) );
  NAND2_X2 U334 ( .A1(n618), .A2(n619), .ZN(n291) );
  NAND2_X1 U335 ( .A1(StartIn), .A2(n811), .ZN(n292) );
  INV_X4 U336 ( .A(n292), .ZN(n293) );
  NAND2_X1 U337 ( .A1(n809), .A2(n814), .ZN(n811) );
  XOR2_X2 U338 ( .A(n298), .B(n354), .Z(n788) );
  INV_X2 U339 ( .A(n783), .ZN(n358) );
  XOR2_X1 U340 ( .A(n610), .B(n759), .Z(n573) );
  NAND2_X2 U341 ( .A1(n619), .A2(n618), .ZN(n735) );
  NAND2_X2 U342 ( .A1(n480), .A2(n295), .ZN(n485) );
  INV_X4 U343 ( .A(n294), .ZN(n295) );
  OR2_X1 U344 ( .A1(n620), .A2(n610), .ZN(n296) );
  NAND4_X4 U345 ( .A1(n421), .A2(n420), .A3(n419), .A4(n418), .ZN(n610) );
  NAND3_X4 U346 ( .A1(n222), .A2(n563), .A3(n221), .ZN(n564) );
  NAND2_X2 U347 ( .A1(n505), .A2(n506), .ZN(n528) );
  NOR2_X2 U348 ( .A1(n330), .A2(n232), .ZN(n300) );
  NAND2_X2 U349 ( .A1(n302), .A2(n301), .ZN(n316) );
  INV_X2 U350 ( .A(CdfMin[0]), .ZN(n375) );
  NAND3_X1 U351 ( .A1(n287), .A2(n402), .A3(n401), .ZN(n458) );
  INV_X2 U352 ( .A(CdfMin[2]), .ZN(n381) );
  NAND2_X2 U353 ( .A1(n539), .A2(n349), .ZN(n311) );
  NAND2_X2 U354 ( .A1(n485), .A2(n486), .ZN(n305) );
  XOR2_X1 U355 ( .A(n252), .B(n351), .Z(n669) );
  XOR2_X1 U356 ( .A(n424), .B(n304), .Z(n410) );
  INV_X1 U357 ( .A(n410), .ZN(n411) );
  NAND3_X1 U358 ( .A1(n527), .A2(n229), .A3(n508), .ZN(n456) );
  NAND2_X2 U359 ( .A1(n542), .A2(n212), .ZN(n488) );
  INV_X4 U360 ( .A(n347), .ZN(n319) );
  INV_X2 U361 ( .A(n713), .ZN(n708) );
  NAND3_X4 U362 ( .A1(n515), .A2(n516), .A3(n517), .ZN(n562) );
  NAND2_X2 U363 ( .A1(n494), .A2(n310), .ZN(n309) );
  NAND3_X2 U364 ( .A1(n312), .A2(n534), .A3(n532), .ZN(n533) );
  INV_X2 U365 ( .A(n311), .ZN(n312) );
  INV_X4 U366 ( .A(n313), .ZN(n314) );
  NAND2_X2 U367 ( .A1(n494), .A2(n310), .ZN(n578) );
  NAND2_X1 U368 ( .A1(n710), .A2(n712), .ZN(n731) );
  NAND2_X2 U369 ( .A1(n374), .A2(DataIn[1]), .ZN(n387) );
  INV_X4 U370 ( .A(CdfMin[1]), .ZN(n374) );
  NAND2_X2 U371 ( .A1(n388), .A2(n387), .ZN(n361) );
  OAI22_X2 U372 ( .A1(n545), .A2(n207), .B1(n614), .B2(n548), .ZN(n566) );
  NOR2_X1 U373 ( .A1(n330), .A2(n583), .ZN(n584) );
  NAND3_X2 U374 ( .A1(n611), .A2(n165), .A3(n612), .ZN(n619) );
  AND2_X1 U375 ( .A1(n783), .A2(n767), .ZN(n317) );
  NOR3_X2 U376 ( .A1(n317), .A2(n318), .A3(n749), .ZN(U4_Z_21) );
  NOR2_X1 U377 ( .A1(n767), .A2(n754), .ZN(n750) );
  INV_X1 U378 ( .A(n594), .ZN(n561) );
  XNOR2_X1 U379 ( .A(CdfMin[14]), .B(DataIn[14]), .ZN(n560) );
  INV_X1 U380 ( .A(n598), .ZN(n559) );
  INV_X1 U381 ( .A(n560), .ZN(n558) );
  XNOR2_X2 U382 ( .A(n305), .B(n319), .ZN(n513) );
  NAND2_X1 U383 ( .A1(n575), .A2(n678), .ZN(n321) );
  NAND2_X2 U384 ( .A1(n320), .A2(n321), .ZN(n612) );
  NAND2_X1 U385 ( .A1(n276), .A2(n452), .ZN(n324) );
  NAND2_X1 U386 ( .A1(n799), .A2(n766), .ZN(n754) );
  OAI221_X2 U387 ( .B1(n652), .B2(n286), .C1(n330), .C2(n232), .A(n651), .ZN(
        n325) );
  AND2_X2 U388 ( .A1(n552), .A2(n577), .ZN(n329) );
  INV_X2 U389 ( .A(n724), .ZN(n332) );
  AND2_X4 U390 ( .A1(n345), .A2(n638), .ZN(n333) );
  AND2_X4 U391 ( .A1(n717), .A2(n719), .ZN(n336) );
  AND2_X4 U392 ( .A1(n206), .A2(n521), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n603), .B(n241), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n231), .B(n789), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n782), .B(n737), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n207), .B(n550), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n713), .B(n650), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n221), .B(n795), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n344), .B(n331), .ZN(n519) );
  XNOR2_X1 U400 ( .A(n289), .B(n482), .ZN(n483) );
  XOR2_X1 U401 ( .A(n708), .B(n226), .Z(n482) );
  XNOR2_X1 U402 ( .A(n476), .B(n737), .ZN(n343) );
  XNOR2_X1 U403 ( .A(CdfMin[16]), .B(DataIn[16]), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n522), .B(CdfMin[11]), .ZN(n354) );
  XNOR2_X1 U405 ( .A(n262), .B(n484), .ZN(n347) );
  OR2_X2 U406 ( .A1(CdfMin[8]), .A2(n348), .ZN(n498) );
  NOR2_X1 U407 ( .A1(n535), .A2(n349), .ZN(n326) );
  NOR2_X1 U408 ( .A1(n534), .A2(n349), .ZN(n327) );
  XNOR2_X1 U409 ( .A(n525), .B(DataIn[12]), .ZN(n349) );
  NAND2_X2 U410 ( .A1(n257), .A2(n766), .ZN(n565) );
  OR3_X1 U411 ( .A1(n715), .A2(n332), .A3(n716), .ZN(n727) );
  INV_X4 U412 ( .A(n366), .ZN(n364) );
  INV_X4 U413 ( .A(n366), .ZN(n365) );
  XNOR2_X2 U414 ( .A(n334), .B(n352), .ZN(n711) );
  XNOR2_X2 U415 ( .A(n335), .B(n660), .ZN(n661) );
  INV_X1 U416 ( .A(n336), .ZN(n668) );
  XNOR2_X2 U417 ( .A(n604), .B(n337), .ZN(n605) );
  XNOR2_X2 U418 ( .A(n338), .B(n806), .ZN(n733) );
  XNOR2_X2 U419 ( .A(n536), .B(n340), .ZN(n537) );
  XNOR2_X2 U420 ( .A(n343), .B(n463), .ZN(n464) );
  AND2_X1 U421 ( .A1(n598), .A2(n597), .ZN(n345) );
  INV_X4 U422 ( .A(reset_n), .ZN(n366) );
  OR2_X1 U423 ( .A1(n683), .A2(CdfMin[18]), .ZN(n690) );
  INV_X4 U424 ( .A(StartIn), .ZN(n804) );
  NAND2_X1 U425 ( .A1(n708), .A2(n709), .ZN(n710) );
  INV_X4 U426 ( .A(n254), .ZN(n357) );
  NAND2_X2 U427 ( .A1(n309), .A2(n579), .ZN(n580) );
  NAND2_X1 U428 ( .A1(n177), .A2(n756), .ZN(n807) );
  NOR3_X2 U429 ( .A1(n771), .A2(n772), .A3(n773), .ZN(n775) );
  NOR2_X1 U430 ( .A1(n759), .A2(n767), .ZN(n751) );
  NOR2_X1 U431 ( .A1(n759), .A2(n768), .ZN(n752) );
  OAI211_X1 U432 ( .C1(n161), .C2(n708), .A(n784), .B(n672), .ZN(n674) );
  NAND3_X1 U433 ( .A1(n673), .A2(n672), .A3(n708), .ZN(n675) );
  OAI21_X1 U434 ( .B1(n708), .B2(n784), .A(n673), .ZN(n670) );
  INV_X1 U435 ( .A(n359), .ZN(n360) );
  NOR2_X2 U436 ( .A1(n225), .A2(n546), .ZN(n545) );
  NAND4_X1 U437 ( .A1(n790), .A2(n789), .A3(n231), .A4(n796), .ZN(n793) );
  NAND3_X1 U438 ( .A1(n741), .A2(n740), .A3(n231), .ZN(n742) );
  XNOR2_X1 U439 ( .A(n495), .B(n204), .ZN(n496) );
  NAND3_X1 U440 ( .A1(n768), .A2(n256), .A3(n767), .ZN(n773) );
  NAND2_X1 U441 ( .A1(n160), .A2(n256), .ZN(n762) );
  NAND2_X2 U442 ( .A1(n387), .A2(n388), .ZN(n446) );
  XOR2_X1 U443 ( .A(n575), .B(n271), .Z(n767) );
  NAND3_X1 U444 ( .A1(n680), .A2(n646), .A3(n271), .ZN(n647) );
  NAND2_X1 U445 ( .A1(n790), .A2(n186), .ZN(n787) );
  NOR2_X1 U446 ( .A1(n524), .A2(n268), .ZN(n535) );
  NAND2_X2 U447 ( .A1(n269), .A2(n732), .ZN(n363) );
  INV_X2 U448 ( .A(n446), .ZN(n389) );
  NAND4_X1 U449 ( .A1(n747), .A2(StartIn), .A3(n768), .A4(n186), .ZN(n745) );
  INV_X1 U450 ( .A(n625), .ZN(n587) );
  NAND2_X1 U451 ( .A1(n333), .A2(n290), .ZN(n679) );
  NAND3_X1 U452 ( .A1(n333), .A2(n644), .A3(n290), .ZN(n649) );
  NAND2_X1 U453 ( .A1(n316), .A2(n387), .ZN(n380) );
  INV_X2 U454 ( .A(n612), .ZN(n576) );
  INV_X4 U455 ( .A(n371), .ZN(U4_Z_0) );
  INV_X4 U456 ( .A(n373), .ZN(n476) );
  NOR2_X2 U457 ( .A1(n370), .A2(n804), .ZN(U4_Z_1) );
  NAND2_X2 U458 ( .A1(n372), .A2(n371), .ZN(n378) );
  INV_X4 U459 ( .A(DataIn[2]), .ZN(n379) );
  OAI22_X2 U460 ( .A1(DataIn[0]), .A2(n375), .B1(n374), .B2(DataIn[1]), .ZN(
        n445) );
  XOR2_X2 U461 ( .A(n469), .B(n376), .Z(n517) );
  MUX2_X2 U462 ( .A(n378), .B(n377), .S(n579), .Z(U4_Z_2) );
  NAND2_X2 U463 ( .A1(n303), .A2(n379), .ZN(n385) );
  NAND2_X2 U464 ( .A1(DataIn[2]), .A2(n381), .ZN(n388) );
  INV_X4 U465 ( .A(n391), .ZN(n405) );
  NOR2_X2 U466 ( .A1(n383), .A2(n804), .ZN(U4_Z_3) );
  INV_X4 U467 ( .A(DataIn[4]), .ZN(n452) );
  NAND2_X2 U468 ( .A1(n385), .A2(n386), .ZN(n399) );
  NAND2_X2 U469 ( .A1(n287), .A2(n202), .ZN(n425) );
  INV_X4 U470 ( .A(CdfMin[3]), .ZN(n390) );
  NAND2_X2 U471 ( .A1(DataIn[3]), .A2(n390), .ZN(n426) );
  XOR2_X2 U472 ( .A(n550), .B(n392), .Z(n393) );
  NOR2_X2 U473 ( .A1(n393), .A2(n804), .ZN(U4_Z_4) );
  INV_X4 U474 ( .A(DataIn[5]), .ZN(n408) );
  INV_X4 U475 ( .A(n396), .ZN(n398) );
  NAND2_X2 U476 ( .A1(DataIn[4]), .A2(n275), .ZN(n441) );
  INV_X4 U477 ( .A(n413), .ZN(n394) );
  NAND2_X2 U478 ( .A1(n442), .A2(n324), .ZN(n395) );
  OAI22_X2 U479 ( .A1(n398), .A2(n397), .B1(n400), .B2(n396), .ZN(n403) );
  NAND3_X2 U480 ( .A1(n404), .A2(n403), .A3(n458), .ZN(n616) );
  INV_X4 U481 ( .A(n616), .ZN(n588) );
  XNOR2_X2 U482 ( .A(n588), .B(n435), .ZN(n406) );
  NOR2_X2 U483 ( .A1(n406), .A2(n804), .ZN(U4_Z_5) );
  INV_X4 U484 ( .A(DataIn[6]), .ZN(n424) );
  NAND2_X2 U485 ( .A1(n453), .A2(n409), .ZN(n412) );
  OAI22_X2 U486 ( .A1(n443), .A2(n411), .B1(n171), .B2(n410), .ZN(n421) );
  NAND2_X2 U487 ( .A1(n416), .A2(n415), .ZN(n417) );
  NAND2_X2 U488 ( .A1(n428), .A2(n468), .ZN(n418) );
  INV_X4 U489 ( .A(n610), .ZN(n461) );
  NOR2_X2 U490 ( .A1(n588), .A2(n435), .ZN(n422) );
  XOR2_X2 U491 ( .A(n461), .B(n422), .Z(n423) );
  NOR2_X2 U492 ( .A1(n423), .A2(n804), .ZN(U4_Z_6) );
  INV_X4 U493 ( .A(n427), .ZN(n434) );
  NAND3_X2 U494 ( .A1(n454), .A2(n426), .A3(n441), .ZN(n429) );
  INV_X4 U495 ( .A(n429), .ZN(n506) );
  OAI33_X1 U496 ( .A1(n433), .A2(n428), .A3(n236), .B1(n427), .B2(n350), .B3(
        n506), .ZN(n430) );
  NOR2_X2 U497 ( .A1(n430), .A2(n431), .ZN(n432) );
  NOR3_X2 U498 ( .A1(n588), .A2(n461), .A3(n435), .ZN(n436) );
  XOR2_X2 U499 ( .A(n241), .B(n436), .Z(n437) );
  NOR2_X2 U500 ( .A1(n437), .A2(n804), .ZN(U4_Z_7) );
  INV_X4 U501 ( .A(n438), .ZN(n439) );
  NAND2_X2 U502 ( .A1(DataIn[7]), .A2(n440), .ZN(n449) );
  OAI21_X4 U503 ( .B1(n447), .B2(n361), .A(n242), .ZN(n505) );
  NAND4_X2 U504 ( .A1(n505), .A2(n448), .A3(n272), .A4(n449), .ZN(n466) );
  NAND2_X2 U505 ( .A1(n457), .A2(n456), .ZN(n465) );
  INV_X4 U506 ( .A(n711), .ZN(n737) );
  INV_X4 U507 ( .A(n458), .ZN(n474) );
  NOR4_X2 U508 ( .A1(n462), .A2(n550), .A3(n241), .A4(n461), .ZN(n463) );
  NOR2_X2 U509 ( .A1(n464), .A2(n804), .ZN(U4_Z_8) );
  NOR4_X2 U510 ( .A1(n472), .A2(n471), .A3(n353), .A4(n350), .ZN(n473) );
  NAND2_X2 U511 ( .A1(n473), .A2(n474), .ZN(n475) );
  NAND2_X2 U512 ( .A1(n475), .A2(n476), .ZN(n489) );
  NAND2_X2 U513 ( .A1(CdfMin[8]), .A2(n348), .ZN(n530) );
  NAND2_X2 U514 ( .A1(n477), .A2(n498), .ZN(n520) );
  INV_X4 U515 ( .A(n520), .ZN(n486) );
  NAND2_X2 U516 ( .A1(n288), .A2(n242), .ZN(n479) );
  NAND2_X2 U517 ( .A1(n479), .A2(n506), .ZN(n480) );
  NOR2_X2 U518 ( .A1(n483), .A2(n804), .ZN(U4_Z_9) );
  NAND2_X2 U519 ( .A1(n486), .A2(n485), .ZN(n542) );
  NAND2_X2 U520 ( .A1(n487), .A2(DataIn[9]), .ZN(n501) );
  INV_X4 U521 ( .A(DataIn[10]), .ZN(n500) );
  INV_X4 U522 ( .A(n512), .ZN(n491) );
  NAND2_X2 U523 ( .A1(n492), .A2(n183), .ZN(n493) );
  NAND2_X2 U524 ( .A1(n493), .A2(n513), .ZN(n494) );
  NOR2_X2 U525 ( .A1(n496), .A2(n804), .ZN(U4_Z_10) );
  NAND2_X2 U526 ( .A1(CdfMin[10]), .A2(n500), .ZN(n499) );
  NAND2_X2 U527 ( .A1(n341), .A2(n530), .ZN(n497) );
  INV_X4 U528 ( .A(DataIn[11]), .ZN(n522) );
  NAND2_X2 U529 ( .A1(n492), .A2(n183), .ZN(n514) );
  XOR2_X2 U530 ( .A(n518), .B(n351), .Z(n721) );
  NOR2_X2 U531 ( .A1(n519), .A2(n804), .ZN(U4_Z_11) );
  NAND2_X2 U532 ( .A1(CdfMin[11]), .A2(n522), .ZN(n521) );
  NAND2_X2 U533 ( .A1(n342), .A2(n520), .ZN(n532) );
  INV_X4 U534 ( .A(n532), .ZN(n524) );
  INV_X4 U535 ( .A(n521), .ZN(n523) );
  OAI22_X2 U536 ( .A1(n248), .A2(n523), .B1(CdfMin[11]), .B2(n522), .ZN(n531)
         );
  INV_X4 U537 ( .A(CdfMin[12]), .ZN(n525) );
  INV_X4 U538 ( .A(n531), .ZN(n539) );
  NOR2_X2 U539 ( .A1(n537), .A2(n804), .ZN(U4_Z_12) );
  INV_X4 U540 ( .A(DataIn[13]), .ZN(n556) );
  XOR2_X2 U541 ( .A(n556), .B(CdfMin[13]), .Z(n575) );
  INV_X4 U542 ( .A(DataIn[12]), .ZN(n538) );
  NAND2_X2 U543 ( .A1(CdfMin[12]), .A2(n538), .ZN(n543) );
  INV_X4 U544 ( .A(n543), .ZN(n540) );
  OAI22_X2 U545 ( .A1(n539), .A2(n540), .B1(CdfMin[12]), .B2(n538), .ZN(n541)
         );
  INV_X4 U546 ( .A(n541), .ZN(n600) );
  INV_X4 U547 ( .A(n767), .ZN(n753) );
  XOR2_X2 U548 ( .A(n616), .B(n753), .Z(n553) );
  XOR2_X2 U549 ( .A(n544), .B(n354), .Z(n547) );
  NAND2_X2 U550 ( .A1(n550), .A2(n788), .ZN(n615) );
  XOR2_X2 U551 ( .A(n553), .B(n329), .Z(n554) );
  NOR2_X2 U552 ( .A1(n554), .A2(n804), .ZN(U4_Z_13) );
  INV_X4 U553 ( .A(CdfMin[13]), .ZN(n555) );
  NAND2_X2 U554 ( .A1(DataIn[13]), .A2(n555), .ZN(n594) );
  NAND2_X2 U555 ( .A1(CdfMin[13]), .A2(n556), .ZN(n598) );
  OAI33_X1 U556 ( .A1(n290), .A2(n561), .A3(n560), .B1(n645), .B2(n559), .B3(
        n558), .ZN(n557) );
  NOR3_X2 U557 ( .A1(n568), .A2(n270), .A3(n567), .ZN(n569) );
  OAI22_X2 U558 ( .A1(n286), .A2(n615), .B1(n570), .B2(n569), .ZN(n611) );
  OAI22_X2 U559 ( .A1(n329), .A2(n616), .B1(n753), .B2(n571), .ZN(n572) );
  INV_X4 U560 ( .A(n572), .ZN(n592) );
  XOR2_X2 U561 ( .A(n592), .B(n573), .Z(n574) );
  NOR2_X2 U562 ( .A1(n574), .A2(n804), .ZN(U4_Z_14) );
  INV_X4 U563 ( .A(n577), .ZN(n585) );
  NOR2_X2 U564 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X2 U565 ( .A1(n588), .A2(n244), .ZN(n589) );
  NAND2_X2 U566 ( .A1(n589), .A2(n610), .ZN(n627) );
  NOR2_X2 U567 ( .A1(n590), .A2(n627), .ZN(n591) );
  INV_X4 U568 ( .A(DataIn[15]), .ZN(n632) );
  XOR2_X2 U569 ( .A(n632), .B(CdfMin[15]), .Z(n607) );
  INV_X4 U570 ( .A(DataIn[14]), .ZN(n593) );
  NAND2_X2 U571 ( .A1(CdfMin[14]), .A2(n593), .ZN(n597) );
  INV_X4 U572 ( .A(n597), .ZN(n595) );
  OAI22_X2 U573 ( .A1(n595), .A2(n594), .B1(CdfMin[14]), .B2(n593), .ZN(n596)
         );
  INV_X4 U574 ( .A(n596), .ZN(n641) );
  NAND2_X2 U575 ( .A1(n641), .A2(n606), .ZN(n633) );
  XOR2_X2 U576 ( .A(n607), .B(n602), .Z(n774) );
  INV_X4 U577 ( .A(n774), .ZN(n603) );
  NOR2_X2 U578 ( .A1(n605), .A2(n804), .ZN(U4_Z_15) );
  NAND2_X2 U579 ( .A1(n281), .A2(n621), .ZN(n623) );
  NAND2_X2 U580 ( .A1(n624), .A2(n625), .ZN(n652) );
  INV_X4 U581 ( .A(n627), .ZN(n629) );
  NAND2_X2 U582 ( .A1(n629), .A2(n628), .ZN(n630) );
  INV_X4 U583 ( .A(n630), .ZN(n651) );
  NAND2_X2 U584 ( .A1(n631), .A2(n308), .ZN(n736) );
  NAND2_X2 U585 ( .A1(CdfMin[15]), .A2(n632), .ZN(n637) );
  INV_X4 U586 ( .A(CdfMin[15]), .ZN(n634) );
  NAND2_X2 U587 ( .A1(DataIn[15]), .A2(n634), .ZN(n701) );
  INV_X4 U588 ( .A(n780), .ZN(n782) );
  NOR2_X2 U589 ( .A1(n635), .A2(n804), .ZN(U4_Z_16) );
  INV_X4 U590 ( .A(DataIn[16]), .ZN(n636) );
  NAND2_X2 U591 ( .A1(CdfMin[16]), .A2(n636), .ZN(n719) );
  NAND2_X2 U592 ( .A1(n719), .A2(n637), .ZN(n640) );
  INV_X4 U593 ( .A(n640), .ZN(n638) );
  INV_X4 U594 ( .A(CdfMin[17]), .ZN(n662) );
  XOR2_X2 U595 ( .A(n662), .B(DataIn[17]), .Z(n644) );
  NOR2_X2 U596 ( .A1(n333), .A2(n644), .ZN(n643) );
  INV_X4 U597 ( .A(n719), .ZN(n723) );
  INV_X4 U598 ( .A(CdfMin[16]), .ZN(n639) );
  NAND2_X2 U599 ( .A1(DataIn[16]), .A2(n639), .ZN(n667) );
  OAI221_X2 U600 ( .B1(n641), .B2(n640), .C1(n723), .C2(n701), .A(n667), .ZN(
        n642) );
  INV_X4 U601 ( .A(n642), .ZN(n680) );
  OAI22_X2 U602 ( .A1(n643), .A2(n642), .B1(n680), .B2(n644), .ZN(n648) );
  INV_X4 U603 ( .A(n644), .ZN(n646) );
  NAND3_X2 U604 ( .A1(n649), .A2(n648), .A3(n647), .ZN(n784) );
  INV_X4 U605 ( .A(n784), .ZN(n650) );
  NAND2_X2 U606 ( .A1(n651), .A2(n737), .ZN(n655) );
  OAI22_X2 U607 ( .A1(n654), .A2(n655), .B1(n308), .B2(n711), .ZN(n656) );
  OAI22_X2 U608 ( .A1(n737), .A2(n659), .B1(n658), .B2(n782), .ZN(n673) );
  NOR2_X2 U609 ( .A1(n661), .A2(n804), .ZN(U4_Z_17) );
  INV_X4 U610 ( .A(DataIn[18]), .ZN(n683) );
  XOR2_X2 U611 ( .A(n683), .B(CdfMin[18]), .Z(n666) );
  INV_X4 U612 ( .A(n666), .ZN(n663) );
  NAND2_X2 U613 ( .A1(DataIn[17]), .A2(n662), .ZN(n685) );
  NAND3_X2 U614 ( .A1(n663), .A2(n667), .A3(n685), .ZN(n724) );
  INV_X4 U615 ( .A(DataIn[17]), .ZN(n664) );
  NAND2_X2 U616 ( .A1(CdfMin[17]), .A2(n664), .ZN(n681) );
  INV_X4 U617 ( .A(n685), .ZN(n691) );
  NAND2_X2 U618 ( .A1(n691), .A2(n666), .ZN(n665) );
  OAI221_X2 U619 ( .B1(n720), .B2(n667), .C1(n666), .C2(n681), .A(n665), .ZN(
        n716) );
  INV_X4 U620 ( .A(n716), .ZN(n722) );
  OAI221_X2 U621 ( .B1(n336), .B2(n724), .C1(n720), .C2(n668), .A(n722), .ZN(
        n796) );
  INV_X4 U622 ( .A(n796), .ZN(n809) );
  XOR2_X2 U623 ( .A(n809), .B(n669), .Z(n672) );
  NAND2_X2 U624 ( .A1(n670), .A2(n671), .ZN(n676) );
  NAND4_X2 U625 ( .A1(n676), .A2(n674), .A3(StartIn), .A4(n675), .ZN(n677) );
  NAND2_X2 U626 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X2 U627 ( .A1(n682), .A2(n681), .ZN(n686) );
  INV_X4 U628 ( .A(n686), .ZN(n684) );
  NAND2_X2 U629 ( .A1(CdfMin[18]), .A2(n683), .ZN(n692) );
  XNOR2_X2 U630 ( .A(CdfMin[19]), .B(DataIn[19]), .ZN(n693) );
  NAND3_X2 U631 ( .A1(n684), .A2(n692), .A3(n693), .ZN(n697) );
  INV_X4 U632 ( .A(n693), .ZN(n687) );
  NAND4_X2 U633 ( .A1(n687), .A2(n686), .A3(n690), .A4(n685), .ZN(n696) );
  INV_X4 U634 ( .A(n690), .ZN(n689) );
  NOR2_X2 U635 ( .A1(n693), .A2(n692), .ZN(n688) );
  OAI22_X2 U636 ( .A1(n693), .A2(n690), .B1(n689), .B2(n688), .ZN(n695) );
  NAND3_X2 U637 ( .A1(n693), .A2(n692), .A3(n691), .ZN(n694) );
  INV_X4 U638 ( .A(n814), .ZN(n789) );
  INV_X4 U639 ( .A(n720), .ZN(n698) );
  NAND2_X2 U640 ( .A1(n698), .A2(n719), .ZN(n703) );
  NOR2_X2 U641 ( .A1(n701), .A2(n703), .ZN(n700) );
  NAND2_X2 U642 ( .A1(n702), .A2(n701), .ZN(n715) );
  NOR2_X2 U643 ( .A1(n724), .A2(n715), .ZN(n705) );
  NAND2_X2 U644 ( .A1(n709), .A2(n784), .ZN(n712) );
  NAND2_X2 U645 ( .A1(n714), .A2(n708), .ZN(n729) );
  INV_X4 U646 ( .A(n716), .ZN(n718) );
  NAND4_X2 U647 ( .A1(n720), .A2(n719), .A3(n718), .A4(n717), .ZN(n726) );
  NAND3_X2 U648 ( .A1(n724), .A2(n723), .A3(n722), .ZN(n725) );
  NAND4_X2 U649 ( .A1(n727), .A2(n726), .A3(n187), .A4(n725), .ZN(n728) );
  NAND2_X2 U650 ( .A1(n736), .A2(n740), .ZN(n730) );
  OAI22_X2 U651 ( .A1(n180), .A2(n739), .B1(n735), .B2(n730), .ZN(n756) );
  INV_X4 U652 ( .A(n741), .ZN(n732) );
  NOR2_X2 U653 ( .A1(n733), .A2(n804), .ZN(U4_Z_19) );
  NOR2_X2 U654 ( .A1(n739), .A2(n795), .ZN(n738) );
  NAND4_X2 U655 ( .A1(n362), .A2(n657), .A3(n738), .A4(n737), .ZN(n743) );
  INV_X4 U656 ( .A(n786), .ZN(n810) );
  NAND2_X2 U657 ( .A1(n207), .A2(StartIn), .ZN(n746) );
  NAND2_X2 U658 ( .A1(n756), .A2(n363), .ZN(n755) );
  NAND2_X2 U659 ( .A1(n795), .A2(n814), .ZN(n799) );
  INV_X4 U660 ( .A(n754), .ZN(n768) );
  NAND2_X2 U661 ( .A1(n807), .A2(n814), .ZN(n747) );
  NAND2_X2 U662 ( .A1(n767), .A2(n814), .ZN(n748) );
  NOR2_X2 U663 ( .A1(n752), .A2(n751), .ZN(n764) );
  NAND2_X2 U664 ( .A1(n755), .A2(n814), .ZN(n770) );
  NAND2_X2 U665 ( .A1(n756), .A2(n363), .ZN(n757) );
  NAND2_X2 U666 ( .A1(n755), .A2(n795), .ZN(n769) );
  NAND4_X2 U667 ( .A1(n763), .A2(StartIn), .A3(n764), .A4(n762), .ZN(n765) );
  NAND4_X2 U668 ( .A1(n774), .A2(n256), .A3(n767), .A4(n766), .ZN(n781) );
  OAI33_X1 U669 ( .A1(n778), .A2(n781), .A3(n804), .B1(n775), .B2(n774), .B3(
        n804), .ZN(n817) );
  NAND2_X2 U670 ( .A1(StartIn), .A2(n776), .ZN(n777) );
  INV_X4 U671 ( .A(n781), .ZN(n779) );
  NAND3_X2 U672 ( .A1(n784), .A2(n780), .A3(n779), .ZN(n815) );
  INV_X4 U673 ( .A(n815), .ZN(n790) );
  NOR4_X2 U674 ( .A1(n357), .A2(n247), .A3(n782), .A4(n781), .ZN(n785) );
  OAI33_X1 U675 ( .A1(n787), .A2(n804), .A3(n159), .B1(n785), .B2(n804), .B3(
        n784), .ZN(n818) );
  INV_X4 U676 ( .A(n811), .ZN(n791) );
  NAND2_X2 U677 ( .A1(n791), .A2(n795), .ZN(n792) );
  NAND2_X2 U678 ( .A1(n793), .A2(n792), .ZN(n803) );
  INV_X4 U679 ( .A(n794), .ZN(n802) );
  NOR2_X2 U680 ( .A1(n795), .A2(n814), .ZN(n797) );
  NOR2_X2 U681 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR3_X2 U682 ( .A1(n803), .A2(n802), .A3(n798), .ZN(n808) );
  INV_X4 U683 ( .A(n799), .ZN(n800) );
  NOR3_X2 U684 ( .A1(n800), .A2(n809), .A3(n815), .ZN(n801) );
  NOR3_X2 U685 ( .A1(n803), .A2(n802), .A3(n801), .ZN(n805) );
  AOI221_X2 U686 ( .B1(n807), .B2(n808), .C1(n806), .C2(n805), .A(n804), .ZN(
        U4_Z_26) );
  AOI221_X2 U687 ( .B1(n815), .B2(n814), .C1(n813), .C2(n358), .A(n812), .ZN(
        U4_Z_27) );
endmodule


module pipleline_stage_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64, n65,
         n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n128, n129, n130, n131, n132, n133, n136, n137, n138, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n157, n158, n160, n161, n162, n163, n164,
         n166, n168, n169, n170, n171, n172, n173, n174, n175, n176, n247,
         n249;

  XNOR2_X2 U3 ( .A(n29), .B(n2), .ZN(SUM[19]) );
  NAND2_X2 U9 ( .A1(n158), .A2(n28), .ZN(n2) );
  NAND2_X2 U12 ( .A1(B[19]), .A2(A[19]), .ZN(n28) );
  XNOR2_X2 U13 ( .A(n36), .B(n3), .ZN(SUM[18]) );
  NAND2_X2 U15 ( .A1(n39), .A2(n32), .ZN(n30) );
  NAND2_X2 U19 ( .A1(n32), .A2(n35), .ZN(n3) );
  NAND2_X2 U22 ( .A1(B[18]), .A2(A[18]), .ZN(n35) );
  XNOR2_X2 U23 ( .A(n43), .B(n4), .ZN(SUM[17]) );
  NAND2_X2 U29 ( .A1(n160), .A2(n42), .ZN(n4) );
  NAND2_X2 U32 ( .A1(B[17]), .A2(A[17]), .ZN(n42) );
  XOR2_X2 U33 ( .A(n5), .B(n1), .Z(SUM[16]) );
  NAND2_X2 U35 ( .A1(n161), .A2(n45), .ZN(n5) );
  NAND2_X2 U38 ( .A1(B[16]), .A2(A[16]), .ZN(n45) );
  XNOR2_X2 U39 ( .A(n55), .B(n6), .ZN(SUM[15]) );
  NAND2_X2 U43 ( .A1(n67), .A2(n51), .ZN(n49) );
  NAND2_X2 U47 ( .A1(n162), .A2(n54), .ZN(n6) );
  NAND2_X2 U50 ( .A1(B[15]), .A2(A[15]), .ZN(n54) );
  XNOR2_X2 U51 ( .A(n64), .B(n7), .ZN(SUM[14]) );
  NAND2_X2 U53 ( .A1(n58), .A2(n85), .ZN(n56) );
  NAND2_X2 U59 ( .A1(n163), .A2(n63), .ZN(n7) );
  NAND2_X2 U62 ( .A1(B[14]), .A2(A[14]), .ZN(n63) );
  XNOR2_X2 U63 ( .A(n75), .B(n8), .ZN(SUM[13]) );
  NAND2_X2 U65 ( .A1(n85), .A2(n67), .ZN(n65) );
  NAND2_X2 U73 ( .A1(n164), .A2(n74), .ZN(n8) );
  NAND2_X2 U76 ( .A1(B[13]), .A2(A[13]), .ZN(n74) );
  XNOR2_X2 U77 ( .A(n82), .B(n9), .ZN(SUM[12]) );
  NAND2_X2 U79 ( .A1(n85), .A2(n78), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n78), .A2(n81), .ZN(n9) );
  NAND2_X2 U86 ( .A1(B[12]), .A2(A[12]), .ZN(n81) );
  XNOR2_X2 U87 ( .A(n93), .B(n10), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(n103), .A2(n89), .ZN(n83) );
  NAND2_X2 U97 ( .A1(n166), .A2(n92), .ZN(n10) );
  NAND2_X2 U100 ( .A1(B[11]), .A2(A[11]), .ZN(n92) );
  XNOR2_X2 U101 ( .A(n100), .B(n11), .ZN(SUM[10]) );
  NAND2_X2 U103 ( .A1(n103), .A2(n96), .ZN(n94) );
  NAND2_X2 U107 ( .A1(n96), .A2(n99), .ZN(n11) );
  NAND2_X2 U110 ( .A1(B[10]), .A2(A[10]), .ZN(n99) );
  XNOR2_X2 U111 ( .A(n111), .B(n12), .ZN(SUM[9]) );
  NAND2_X2 U121 ( .A1(n168), .A2(n110), .ZN(n12) );
  NAND2_X2 U124 ( .A1(B[9]), .A2(A[9]), .ZN(n110) );
  XOR2_X2 U125 ( .A(n13), .B(n114), .Z(SUM[8]) );
  NAND2_X2 U127 ( .A1(n169), .A2(n113), .ZN(n13) );
  NAND2_X2 U130 ( .A1(B[8]), .A2(A[8]), .ZN(n113) );
  XOR2_X2 U131 ( .A(n14), .B(n122), .Z(SUM[7]) );
  NAND2_X2 U134 ( .A1(n130), .A2(n118), .ZN(n116) );
  NAND2_X2 U138 ( .A1(n170), .A2(n121), .ZN(n14) );
  NAND2_X2 U141 ( .A1(B[7]), .A2(A[7]), .ZN(n121) );
  XOR2_X2 U142 ( .A(n15), .B(n129), .Z(SUM[6]) );
  NAND2_X2 U148 ( .A1(n171), .A2(n128), .ZN(n15) );
  NAND2_X2 U151 ( .A1(B[6]), .A2(A[6]), .ZN(n128) );
  XOR2_X2 U152 ( .A(n16), .B(n138), .Z(SUM[5]) );
  NAND2_X2 U160 ( .A1(n172), .A2(n137), .ZN(n16) );
  NAND2_X2 U163 ( .A1(B[5]), .A2(A[5]), .ZN(n137) );
  XNOR2_X2 U164 ( .A(n143), .B(n17), .ZN(SUM[4]) );
  NAND2_X2 U168 ( .A1(n173), .A2(n142), .ZN(n17) );
  NAND2_X2 U171 ( .A1(B[4]), .A2(A[4]), .ZN(n142) );
  XNOR2_X2 U172 ( .A(n149), .B(n18), .ZN(SUM[3]) );
  NAND2_X2 U177 ( .A1(n174), .A2(n148), .ZN(n18) );
  NAND2_X2 U180 ( .A1(B[3]), .A2(A[3]), .ZN(n148) );
  XOR2_X2 U181 ( .A(n19), .B(n152), .Z(SUM[2]) );
  NAND2_X2 U183 ( .A1(n175), .A2(n151), .ZN(n19) );
  NAND2_X2 U186 ( .A1(B[2]), .A2(A[2]), .ZN(n151) );
  XOR2_X2 U187 ( .A(n157), .B(n20), .Z(SUM[1]) );
  NAND2_X2 U190 ( .A1(n176), .A2(n155), .ZN(n20) );
  NAND2_X2 U193 ( .A1(B[1]), .A2(A[1]), .ZN(n155) );
  NAND2_X2 U198 ( .A1(B[0]), .A2(A[0]), .ZN(n157) );
  OR2_X1 U202 ( .A1(n30), .A2(n27), .ZN(n247) );
  AND2_X1 U203 ( .A1(n249), .A2(n157), .ZN(SUM[0]) );
  NOR2_X1 U204 ( .A1(B[2]), .A2(A[2]), .ZN(n150) );
  OAI21_X1 U205 ( .B1(n1), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U206 ( .B1(n114), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X1 U207 ( .B1(n86), .B2(n78), .A(n79), .ZN(n77) );
  AOI21_X1 U208 ( .B1(n86), .B2(n67), .A(n68), .ZN(n66) );
  INV_X1 U209 ( .A(n104), .ZN(n102) );
  AOI21_X1 U210 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  INV_X1 U211 ( .A(n40), .ZN(n38) );
  AOI21_X4 U212 ( .B1(n115), .B2(n47), .A(n48), .ZN(n1) );
  NOR2_X1 U213 ( .A1(n83), .A2(n49), .ZN(n47) );
  NOR2_X1 U214 ( .A1(n150), .A2(n147), .ZN(n145) );
  OAI21_X1 U215 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  OAI21_X1 U216 ( .B1(n133), .B2(n125), .A(n128), .ZN(n124) );
  AOI21_X1 U217 ( .B1(n143), .B2(n123), .A(n124), .ZN(n122) );
  NOR2_X1 U218 ( .A1(n132), .A2(n125), .ZN(n123) );
  NOR2_X1 U219 ( .A1(n80), .A2(n73), .ZN(n67) );
  OAI21_X1 U220 ( .B1(n1), .B2(n44), .A(n45), .ZN(n43) );
  NOR2_X1 U221 ( .A1(n69), .A2(n60), .ZN(n58) );
  OAI21_X1 U222 ( .B1(n114), .B2(n56), .A(n57), .ZN(n55) );
  OAI21_X1 U223 ( .B1(n114), .B2(n94), .A(n95), .ZN(n93) );
  NOR2_X1 U224 ( .A1(n141), .A2(n136), .ZN(n130) );
  NOR2_X1 U225 ( .A1(n112), .A2(n109), .ZN(n103) );
  OAI21_X1 U226 ( .B1(n120), .B2(n128), .A(n121), .ZN(n119) );
  NOR2_X1 U227 ( .A1(n44), .A2(n41), .ZN(n39) );
  NOR2_X1 U228 ( .A1(n98), .A2(n91), .ZN(n89) );
  NOR2_X1 U229 ( .A1(n60), .A2(n53), .ZN(n51) );
  OAI21_X1 U230 ( .B1(n31), .B2(n27), .A(n28), .ZN(n26) );
  NOR2_X1 U231 ( .A1(B[16]), .A2(A[16]), .ZN(n44) );
  NOR2_X1 U232 ( .A1(B[12]), .A2(A[12]), .ZN(n80) );
  OAI21_X2 U233 ( .B1(n84), .B2(n49), .A(n50), .ZN(n48) );
  OAI21_X1 U234 ( .B1(n114), .B2(n101), .A(n102), .ZN(n100) );
  OAI21_X1 U235 ( .B1(n1), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X1 U236 ( .B1(n114), .B2(n83), .A(n84), .ZN(n82) );
  OAI21_X1 U237 ( .B1(n114), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X2 U238 ( .B1(n89), .B2(n104), .A(n90), .ZN(n84) );
  OAI21_X2 U239 ( .B1(n91), .B2(n99), .A(n92), .ZN(n90) );
  AOI21_X1 U240 ( .B1(n40), .B2(n32), .A(n33), .ZN(n31) );
  OAI21_X2 U241 ( .B1(n109), .B2(n113), .A(n110), .ZN(n104) );
  AOI21_X2 U242 ( .B1(n145), .B2(n153), .A(n146), .ZN(n144) );
  OAI21_X2 U243 ( .B1(n73), .B2(n81), .A(n74), .ZN(n68) );
  OAI21_X2 U244 ( .B1(n136), .B2(n142), .A(n137), .ZN(n131) );
  OAI21_X2 U245 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI21_X2 U246 ( .B1(n144), .B2(n116), .A(n117), .ZN(n115) );
  AOI21_X2 U247 ( .B1(n118), .B2(n131), .A(n119), .ZN(n117) );
  NOR2_X2 U248 ( .A1(n125), .A2(n120), .ZN(n118) );
  AOI21_X2 U249 ( .B1(n51), .B2(n68), .A(n52), .ZN(n50) );
  OAI21_X2 U250 ( .B1(n53), .B2(n63), .A(n54), .ZN(n52) );
  AOI21_X2 U251 ( .B1(n143), .B2(n173), .A(n140), .ZN(n138) );
  OAI21_X2 U252 ( .B1(n154), .B2(n157), .A(n155), .ZN(n153) );
  OAI21_X1 U253 ( .B1(n70), .B2(n60), .A(n63), .ZN(n59) );
  OAI21_X1 U254 ( .B1(n114), .B2(n112), .A(n113), .ZN(n111) );
  AOI21_X2 U255 ( .B1(n86), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X1 U256 ( .B1(n104), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U257 ( .B1(n152), .B2(n150), .A(n151), .ZN(n149) );
  NOR2_X2 U258 ( .A1(B[14]), .A2(A[14]), .ZN(n60) );
  NOR2_X2 U259 ( .A1(B[6]), .A2(A[6]), .ZN(n125) );
  NOR2_X2 U260 ( .A1(B[5]), .A2(A[5]), .ZN(n136) );
  NOR2_X2 U261 ( .A1(B[7]), .A2(A[7]), .ZN(n120) );
  NOR2_X2 U262 ( .A1(B[3]), .A2(A[3]), .ZN(n147) );
  NOR2_X2 U263 ( .A1(B[13]), .A2(A[13]), .ZN(n73) );
  NOR2_X2 U264 ( .A1(B[11]), .A2(A[11]), .ZN(n91) );
  NOR2_X2 U265 ( .A1(B[15]), .A2(A[15]), .ZN(n53) );
  NOR2_X2 U266 ( .A1(B[9]), .A2(A[9]), .ZN(n109) );
  NOR2_X2 U267 ( .A1(B[17]), .A2(A[17]), .ZN(n41) );
  NOR2_X2 U268 ( .A1(B[19]), .A2(A[19]), .ZN(n27) );
  NOR2_X1 U269 ( .A1(B[8]), .A2(A[8]), .ZN(n112) );
  NOR2_X2 U270 ( .A1(B[1]), .A2(A[1]), .ZN(n154) );
  NOR2_X1 U271 ( .A1(B[4]), .A2(A[4]), .ZN(n141) );
  NOR2_X1 U272 ( .A1(B[10]), .A2(A[10]), .ZN(n98) );
  OAI21_X2 U273 ( .B1(n1), .B2(n247), .A(n24), .ZN(SUM[20]) );
  NOR2_X2 U274 ( .A1(B[18]), .A2(A[18]), .ZN(n34) );
  OR2_X1 U275 ( .A1(B[0]), .A2(A[0]), .ZN(n249) );
  INV_X4 U276 ( .A(n99), .ZN(n97) );
  INV_X4 U277 ( .A(n84), .ZN(n86) );
  INV_X4 U278 ( .A(n83), .ZN(n85) );
  INV_X4 U279 ( .A(n81), .ZN(n79) );
  INV_X4 U280 ( .A(n68), .ZN(n70) );
  INV_X4 U281 ( .A(n67), .ZN(n69) );
  INV_X4 U282 ( .A(n39), .ZN(n37) );
  INV_X4 U283 ( .A(n35), .ZN(n33) );
  INV_X4 U284 ( .A(n26), .ZN(n24) );
  INV_X4 U285 ( .A(n154), .ZN(n176) );
  INV_X4 U286 ( .A(n150), .ZN(n175) );
  INV_X4 U287 ( .A(n147), .ZN(n174) );
  INV_X4 U288 ( .A(n136), .ZN(n172) );
  INV_X4 U289 ( .A(n125), .ZN(n171) );
  INV_X4 U290 ( .A(n120), .ZN(n170) );
  INV_X4 U291 ( .A(n112), .ZN(n169) );
  INV_X4 U292 ( .A(n109), .ZN(n168) );
  INV_X4 U293 ( .A(n98), .ZN(n96) );
  INV_X4 U294 ( .A(n91), .ZN(n166) );
  INV_X4 U295 ( .A(n80), .ZN(n78) );
  INV_X4 U296 ( .A(n73), .ZN(n164) );
  INV_X4 U297 ( .A(n60), .ZN(n163) );
  INV_X4 U298 ( .A(n53), .ZN(n162) );
  INV_X4 U299 ( .A(n44), .ZN(n161) );
  INV_X4 U300 ( .A(n41), .ZN(n160) );
  INV_X4 U301 ( .A(n34), .ZN(n32) );
  INV_X4 U302 ( .A(n27), .ZN(n158) );
  INV_X4 U303 ( .A(n153), .ZN(n152) );
  INV_X4 U304 ( .A(n144), .ZN(n143) );
  INV_X4 U305 ( .A(n142), .ZN(n140) );
  INV_X4 U306 ( .A(n141), .ZN(n173) );
  INV_X4 U307 ( .A(n131), .ZN(n133) );
  INV_X4 U308 ( .A(n130), .ZN(n132) );
  INV_X4 U309 ( .A(n115), .ZN(n114) );
  INV_X4 U310 ( .A(n103), .ZN(n101) );
endmodule


module pipleline_stage_1 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n106;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;

  pipleline_stage_1_DW01_add_1 add_268 ( .A({1'b0, divided[26:7]}), .B({1'b0, 
        divisor}), .CI(1'b0), .SUM(stage_result) );
  BUF_X4 U5 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U6 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U7 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U8 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U9 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U10 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U11 ( .A(divided[0]), .Z(stage_out[1]) );
  INV_X16 U12 ( .A(n106), .ZN(q) );
  XNOR2_X2 U13 ( .A(divided[27]), .B(stage_result[20]), .ZN(n106) );
  MUX2_X2 U14 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U15 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U16 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U17 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U18 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U19 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U20 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U21 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U22 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U23 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U24 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U25 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U26 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U27 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U28 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U29 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U30 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U31 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U32 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U33 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_7_DW01_add_1 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n24, n26, n27, n28, n29, n30, n31, n33, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64, n65, n66, n67,
         n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n128, n129, n130, n131, n132, n133, n136, n137, n138, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n157, n158, n160, n161, n162, n163, n164, n166,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n247, n249,
         n250;

  XNOR2_X2 U3 ( .A(n29), .B(n2), .ZN(SUM[19]) );
  NAND2_X2 U9 ( .A1(n158), .A2(n28), .ZN(n2) );
  NAND2_X2 U12 ( .A1(A[19]), .A2(B[19]), .ZN(n28) );
  XNOR2_X2 U13 ( .A(n36), .B(n3), .ZN(SUM[18]) );
  NAND2_X2 U15 ( .A1(n39), .A2(n249), .ZN(n30) );
  NAND2_X2 U19 ( .A1(n249), .A2(n35), .ZN(n3) );
  NAND2_X2 U22 ( .A1(A[18]), .A2(B[18]), .ZN(n35) );
  XNOR2_X2 U23 ( .A(n43), .B(n4), .ZN(SUM[17]) );
  NAND2_X2 U29 ( .A1(n160), .A2(n42), .ZN(n4) );
  NAND2_X2 U32 ( .A1(A[17]), .A2(B[17]), .ZN(n42) );
  XOR2_X2 U33 ( .A(n5), .B(n1), .Z(SUM[16]) );
  NAND2_X2 U35 ( .A1(n161), .A2(n45), .ZN(n5) );
  NAND2_X2 U38 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U39 ( .A(n55), .B(n6), .ZN(SUM[15]) );
  NAND2_X2 U43 ( .A1(n67), .A2(n51), .ZN(n49) );
  NAND2_X2 U47 ( .A1(n162), .A2(n54), .ZN(n6) );
  NAND2_X2 U50 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  XNOR2_X2 U51 ( .A(n64), .B(n7), .ZN(SUM[14]) );
  NAND2_X2 U53 ( .A1(n58), .A2(n85), .ZN(n56) );
  NAND2_X2 U59 ( .A1(n163), .A2(n63), .ZN(n7) );
  NAND2_X2 U62 ( .A1(A[14]), .A2(B[14]), .ZN(n63) );
  XNOR2_X2 U63 ( .A(n75), .B(n8), .ZN(SUM[13]) );
  NAND2_X2 U65 ( .A1(n85), .A2(n67), .ZN(n65) );
  NAND2_X2 U73 ( .A1(n164), .A2(n74), .ZN(n8) );
  NAND2_X2 U76 ( .A1(A[13]), .A2(B[13]), .ZN(n74) );
  XNOR2_X2 U77 ( .A(n82), .B(n9), .ZN(SUM[12]) );
  NAND2_X2 U79 ( .A1(n85), .A2(n78), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n78), .A2(n81), .ZN(n9) );
  NAND2_X2 U86 ( .A1(A[12]), .A2(B[12]), .ZN(n81) );
  XNOR2_X2 U87 ( .A(n93), .B(n10), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(n103), .A2(n89), .ZN(n83) );
  NAND2_X2 U97 ( .A1(n166), .A2(n92), .ZN(n10) );
  NAND2_X2 U100 ( .A1(A[11]), .A2(B[11]), .ZN(n92) );
  XNOR2_X2 U101 ( .A(n100), .B(n11), .ZN(SUM[10]) );
  NAND2_X2 U103 ( .A1(n103), .A2(n96), .ZN(n94) );
  NAND2_X2 U107 ( .A1(n96), .A2(n99), .ZN(n11) );
  NAND2_X2 U110 ( .A1(A[10]), .A2(B[10]), .ZN(n99) );
  XNOR2_X2 U111 ( .A(n111), .B(n12), .ZN(SUM[9]) );
  NAND2_X2 U121 ( .A1(n168), .A2(n110), .ZN(n12) );
  NAND2_X2 U124 ( .A1(A[9]), .A2(B[9]), .ZN(n110) );
  XOR2_X2 U125 ( .A(n13), .B(n114), .Z(SUM[8]) );
  NAND2_X2 U127 ( .A1(n169), .A2(n113), .ZN(n13) );
  NAND2_X2 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n113) );
  XOR2_X2 U131 ( .A(n14), .B(n122), .Z(SUM[7]) );
  NAND2_X2 U134 ( .A1(n130), .A2(n118), .ZN(n116) );
  NAND2_X2 U138 ( .A1(n170), .A2(n121), .ZN(n14) );
  NAND2_X2 U141 ( .A1(A[7]), .A2(B[7]), .ZN(n121) );
  XOR2_X2 U142 ( .A(n15), .B(n129), .Z(SUM[6]) );
  NAND2_X2 U148 ( .A1(n171), .A2(n128), .ZN(n15) );
  NAND2_X2 U151 ( .A1(A[6]), .A2(B[6]), .ZN(n128) );
  XOR2_X2 U152 ( .A(n16), .B(n138), .Z(SUM[5]) );
  NAND2_X2 U160 ( .A1(n172), .A2(n137), .ZN(n16) );
  NAND2_X2 U163 ( .A1(A[5]), .A2(B[5]), .ZN(n137) );
  XNOR2_X2 U164 ( .A(n143), .B(n17), .ZN(SUM[4]) );
  NAND2_X2 U168 ( .A1(n173), .A2(n142), .ZN(n17) );
  NAND2_X2 U171 ( .A1(A[4]), .A2(B[4]), .ZN(n142) );
  XNOR2_X2 U172 ( .A(n149), .B(n18), .ZN(SUM[3]) );
  NAND2_X2 U177 ( .A1(n174), .A2(n148), .ZN(n18) );
  NAND2_X2 U180 ( .A1(A[3]), .A2(B[3]), .ZN(n148) );
  XOR2_X2 U181 ( .A(n19), .B(n152), .Z(SUM[2]) );
  NAND2_X2 U183 ( .A1(n175), .A2(n151), .ZN(n19) );
  NAND2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n151) );
  XOR2_X2 U187 ( .A(n157), .B(n20), .Z(SUM[1]) );
  NAND2_X2 U190 ( .A1(n176), .A2(n155), .ZN(n20) );
  NAND2_X2 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n155) );
  NAND2_X2 U198 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  OR2_X4 U202 ( .A1(n30), .A2(n27), .ZN(n247) );
  AND2_X1 U203 ( .A1(n250), .A2(n157), .ZN(SUM[0]) );
  NOR2_X1 U204 ( .A1(A[16]), .A2(B[16]), .ZN(n44) );
  NOR2_X1 U205 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  OAI21_X1 U206 ( .B1(n114), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X1 U207 ( .B1(n86), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U208 ( .B1(n114), .B2(n56), .A(n57), .ZN(n55) );
  NOR2_X1 U209 ( .A1(n69), .A2(n60), .ZN(n58) );
  AOI21_X4 U210 ( .B1(n115), .B2(n47), .A(n48), .ZN(n1) );
  NOR2_X1 U211 ( .A1(n83), .A2(n49), .ZN(n47) );
  AOI21_X1 U212 ( .B1(n86), .B2(n67), .A(n68), .ZN(n66) );
  AOI21_X1 U213 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U214 ( .B1(n1), .B2(n37), .A(n38), .ZN(n36) );
  INV_X1 U215 ( .A(n40), .ZN(n38) );
  OAI21_X1 U216 ( .B1(n114), .B2(n101), .A(n102), .ZN(n100) );
  INV_X1 U217 ( .A(n104), .ZN(n102) );
  NOR2_X1 U218 ( .A1(n150), .A2(n147), .ZN(n145) );
  OAI21_X1 U219 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  OAI21_X1 U220 ( .B1(n133), .B2(n125), .A(n128), .ZN(n124) );
  NOR2_X1 U221 ( .A1(n132), .A2(n125), .ZN(n123) );
  NOR2_X1 U222 ( .A1(n80), .A2(n73), .ZN(n67) );
  OAI21_X1 U223 ( .B1(n114), .B2(n94), .A(n95), .ZN(n93) );
  OAI21_X1 U224 ( .B1(n1), .B2(n44), .A(n45), .ZN(n43) );
  NOR2_X1 U225 ( .A1(n141), .A2(n136), .ZN(n130) );
  NOR2_X1 U226 ( .A1(n112), .A2(n109), .ZN(n103) );
  OAI21_X1 U227 ( .B1(n120), .B2(n128), .A(n121), .ZN(n119) );
  NOR2_X1 U228 ( .A1(n44), .A2(n41), .ZN(n39) );
  NOR2_X1 U229 ( .A1(n98), .A2(n91), .ZN(n89) );
  NOR2_X1 U230 ( .A1(n60), .A2(n53), .ZN(n51) );
  OR2_X2 U231 ( .A1(A[18]), .A2(B[18]), .ZN(n249) );
  OAI21_X2 U232 ( .B1(n84), .B2(n49), .A(n50), .ZN(n48) );
  OAI21_X1 U233 ( .B1(n1), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X1 U234 ( .B1(n114), .B2(n83), .A(n84), .ZN(n82) );
  OAI21_X1 U235 ( .B1(n114), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X2 U236 ( .B1(n40), .B2(n249), .A(n33), .ZN(n31) );
  OAI21_X2 U237 ( .B1(n109), .B2(n113), .A(n110), .ZN(n104) );
  AOI21_X2 U238 ( .B1(n145), .B2(n153), .A(n146), .ZN(n144) );
  OAI21_X2 U239 ( .B1(n73), .B2(n81), .A(n74), .ZN(n68) );
  OAI21_X2 U240 ( .B1(n136), .B2(n142), .A(n137), .ZN(n131) );
  OAI21_X2 U241 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI21_X2 U242 ( .B1(n144), .B2(n116), .A(n117), .ZN(n115) );
  AOI21_X2 U243 ( .B1(n118), .B2(n131), .A(n119), .ZN(n117) );
  NOR2_X2 U244 ( .A1(n125), .A2(n120), .ZN(n118) );
  AOI21_X2 U245 ( .B1(n51), .B2(n68), .A(n52), .ZN(n50) );
  OAI21_X2 U246 ( .B1(n53), .B2(n63), .A(n54), .ZN(n52) );
  AOI21_X2 U247 ( .B1(n143), .B2(n123), .A(n124), .ZN(n122) );
  AOI21_X2 U248 ( .B1(n143), .B2(n173), .A(n140), .ZN(n138) );
  OAI21_X2 U249 ( .B1(n154), .B2(n157), .A(n155), .ZN(n153) );
  AOI21_X2 U250 ( .B1(n89), .B2(n104), .A(n90), .ZN(n84) );
  OAI21_X2 U251 ( .B1(n91), .B2(n99), .A(n92), .ZN(n90) );
  OAI21_X1 U252 ( .B1(n70), .B2(n60), .A(n63), .ZN(n59) );
  AOI21_X2 U253 ( .B1(n86), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X1 U254 ( .B1(n104), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U255 ( .B1(n114), .B2(n112), .A(n113), .ZN(n111) );
  OAI21_X1 U256 ( .B1(n152), .B2(n150), .A(n151), .ZN(n149) );
  OAI21_X2 U257 ( .B1(n31), .B2(n27), .A(n28), .ZN(n26) );
  NOR2_X2 U258 ( .A1(A[14]), .A2(B[14]), .ZN(n60) );
  NOR2_X2 U259 ( .A1(A[6]), .A2(B[6]), .ZN(n125) );
  NOR2_X2 U260 ( .A1(A[13]), .A2(B[13]), .ZN(n73) );
  NOR2_X2 U261 ( .A1(A[11]), .A2(B[11]), .ZN(n91) );
  NOR2_X2 U262 ( .A1(A[15]), .A2(B[15]), .ZN(n53) );
  NOR2_X2 U263 ( .A1(A[9]), .A2(B[9]), .ZN(n109) );
  NOR2_X2 U264 ( .A1(A[5]), .A2(B[5]), .ZN(n136) );
  NOR2_X2 U265 ( .A1(A[7]), .A2(B[7]), .ZN(n120) );
  NOR2_X2 U266 ( .A1(A[17]), .A2(B[17]), .ZN(n41) );
  NOR2_X2 U267 ( .A1(A[3]), .A2(B[3]), .ZN(n147) );
  NOR2_X2 U268 ( .A1(A[19]), .A2(B[19]), .ZN(n27) );
  NOR2_X1 U269 ( .A1(A[8]), .A2(B[8]), .ZN(n112) );
  NOR2_X2 U270 ( .A1(A[1]), .A2(B[1]), .ZN(n154) );
  NOR2_X1 U271 ( .A1(A[12]), .A2(B[12]), .ZN(n80) );
  NOR2_X1 U272 ( .A1(A[10]), .A2(B[10]), .ZN(n98) );
  NOR2_X1 U273 ( .A1(A[4]), .A2(B[4]), .ZN(n141) );
  OAI21_X2 U274 ( .B1(n1), .B2(n247), .A(n24), .ZN(SUM[20]) );
  OR2_X1 U275 ( .A1(A[0]), .A2(B[0]), .ZN(n250) );
  INV_X4 U276 ( .A(n99), .ZN(n97) );
  INV_X4 U277 ( .A(n84), .ZN(n86) );
  INV_X4 U278 ( .A(n83), .ZN(n85) );
  INV_X4 U279 ( .A(n81), .ZN(n79) );
  INV_X4 U280 ( .A(n68), .ZN(n70) );
  INV_X4 U281 ( .A(n67), .ZN(n69) );
  INV_X4 U282 ( .A(n39), .ZN(n37) );
  INV_X4 U283 ( .A(n35), .ZN(n33) );
  INV_X4 U284 ( .A(n26), .ZN(n24) );
  INV_X4 U285 ( .A(n154), .ZN(n176) );
  INV_X4 U286 ( .A(n150), .ZN(n175) );
  INV_X4 U287 ( .A(n147), .ZN(n174) );
  INV_X4 U288 ( .A(n136), .ZN(n172) );
  INV_X4 U289 ( .A(n125), .ZN(n171) );
  INV_X4 U290 ( .A(n120), .ZN(n170) );
  INV_X4 U291 ( .A(n112), .ZN(n169) );
  INV_X4 U292 ( .A(n109), .ZN(n168) );
  INV_X4 U293 ( .A(n98), .ZN(n96) );
  INV_X4 U294 ( .A(n91), .ZN(n166) );
  INV_X4 U295 ( .A(n80), .ZN(n78) );
  INV_X4 U296 ( .A(n73), .ZN(n164) );
  INV_X4 U297 ( .A(n60), .ZN(n163) );
  INV_X4 U298 ( .A(n53), .ZN(n162) );
  INV_X4 U299 ( .A(n44), .ZN(n161) );
  INV_X4 U300 ( .A(n41), .ZN(n160) );
  INV_X4 U301 ( .A(n27), .ZN(n158) );
  INV_X4 U302 ( .A(n153), .ZN(n152) );
  INV_X4 U303 ( .A(n144), .ZN(n143) );
  INV_X4 U304 ( .A(n142), .ZN(n140) );
  INV_X4 U305 ( .A(n141), .ZN(n173) );
  INV_X4 U306 ( .A(n131), .ZN(n133) );
  INV_X4 U307 ( .A(n130), .ZN(n132) );
  INV_X4 U308 ( .A(n115), .ZN(n114) );
  INV_X4 U309 ( .A(n103), .ZN(n101) );
endmodule


module pipleline_stage_7 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n106;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;

  pipleline_stage_7_DW01_add_1 add_268 ( .A({1'b0, divided[26:7]}), .B({1'b0, 
        divisor}), .CI(1'b0), .SUM(stage_result) );
  BUF_X4 U5 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U6 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U7 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U8 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U9 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U10 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U11 ( .A(divided[0]), .Z(stage_out[1]) );
  INV_X16 U12 ( .A(n106), .ZN(q) );
  XNOR2_X2 U13 ( .A(divided[27]), .B(stage_result[20]), .ZN(n106) );
  MUX2_X2 U14 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U15 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U16 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U17 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U18 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U19 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U20 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U21 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U22 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U23 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U24 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U25 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U26 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U27 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U28 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U29 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U30 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U31 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U32 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U33 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_6_DW01_add_1 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n24, n26, n27, n28, n29, n30, n31, n33, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64, n65, n66, n67,
         n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n128, n129, n130, n131, n132, n133, n136, n137, n138, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n157, n158, n160, n161, n162, n163, n164, n166,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n247, n248,
         n250;

  XNOR2_X2 U3 ( .A(n29), .B(n2), .ZN(SUM[19]) );
  NAND2_X2 U9 ( .A1(n158), .A2(n28), .ZN(n2) );
  NAND2_X2 U12 ( .A1(A[19]), .A2(B[19]), .ZN(n28) );
  XNOR2_X2 U13 ( .A(n36), .B(n3), .ZN(SUM[18]) );
  NAND2_X2 U15 ( .A1(n39), .A2(n247), .ZN(n30) );
  NAND2_X2 U19 ( .A1(n247), .A2(n35), .ZN(n3) );
  NAND2_X2 U22 ( .A1(A[18]), .A2(B[18]), .ZN(n35) );
  XNOR2_X2 U23 ( .A(n43), .B(n4), .ZN(SUM[17]) );
  NAND2_X2 U29 ( .A1(n160), .A2(n42), .ZN(n4) );
  NAND2_X2 U32 ( .A1(A[17]), .A2(B[17]), .ZN(n42) );
  XOR2_X2 U33 ( .A(n5), .B(n1), .Z(SUM[16]) );
  NAND2_X2 U35 ( .A1(n161), .A2(n45), .ZN(n5) );
  NAND2_X2 U38 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U39 ( .A(n55), .B(n6), .ZN(SUM[15]) );
  NAND2_X2 U43 ( .A1(n67), .A2(n51), .ZN(n49) );
  NAND2_X2 U47 ( .A1(n162), .A2(n54), .ZN(n6) );
  NAND2_X2 U50 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  XNOR2_X2 U51 ( .A(n64), .B(n7), .ZN(SUM[14]) );
  NAND2_X2 U53 ( .A1(n58), .A2(n85), .ZN(n56) );
  NAND2_X2 U59 ( .A1(n163), .A2(n63), .ZN(n7) );
  NAND2_X2 U62 ( .A1(A[14]), .A2(B[14]), .ZN(n63) );
  XNOR2_X2 U63 ( .A(n75), .B(n8), .ZN(SUM[13]) );
  NAND2_X2 U65 ( .A1(n85), .A2(n67), .ZN(n65) );
  NAND2_X2 U73 ( .A1(n164), .A2(n74), .ZN(n8) );
  NAND2_X2 U76 ( .A1(A[13]), .A2(B[13]), .ZN(n74) );
  XNOR2_X2 U77 ( .A(n82), .B(n9), .ZN(SUM[12]) );
  NAND2_X2 U79 ( .A1(n85), .A2(n78), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n78), .A2(n81), .ZN(n9) );
  NAND2_X2 U86 ( .A1(A[12]), .A2(B[12]), .ZN(n81) );
  XNOR2_X2 U87 ( .A(n93), .B(n10), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(n103), .A2(n89), .ZN(n83) );
  NAND2_X2 U97 ( .A1(n166), .A2(n92), .ZN(n10) );
  NAND2_X2 U100 ( .A1(A[11]), .A2(B[11]), .ZN(n92) );
  XNOR2_X2 U101 ( .A(n100), .B(n11), .ZN(SUM[10]) );
  NAND2_X2 U103 ( .A1(n103), .A2(n96), .ZN(n94) );
  NAND2_X2 U107 ( .A1(n96), .A2(n99), .ZN(n11) );
  NAND2_X2 U110 ( .A1(A[10]), .A2(B[10]), .ZN(n99) );
  XNOR2_X2 U111 ( .A(n111), .B(n12), .ZN(SUM[9]) );
  NAND2_X2 U121 ( .A1(n168), .A2(n110), .ZN(n12) );
  NAND2_X2 U124 ( .A1(A[9]), .A2(B[9]), .ZN(n110) );
  XOR2_X2 U125 ( .A(n13), .B(n114), .Z(SUM[8]) );
  NAND2_X2 U127 ( .A1(n169), .A2(n113), .ZN(n13) );
  NAND2_X2 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n113) );
  XOR2_X2 U131 ( .A(n14), .B(n122), .Z(SUM[7]) );
  NAND2_X2 U134 ( .A1(n130), .A2(n118), .ZN(n116) );
  NAND2_X2 U138 ( .A1(n170), .A2(n121), .ZN(n14) );
  NAND2_X2 U141 ( .A1(A[7]), .A2(B[7]), .ZN(n121) );
  XOR2_X2 U142 ( .A(n15), .B(n129), .Z(SUM[6]) );
  NAND2_X2 U148 ( .A1(n171), .A2(n128), .ZN(n15) );
  NAND2_X2 U151 ( .A1(A[6]), .A2(B[6]), .ZN(n128) );
  XOR2_X2 U152 ( .A(n16), .B(n138), .Z(SUM[5]) );
  NAND2_X2 U160 ( .A1(n172), .A2(n137), .ZN(n16) );
  NAND2_X2 U163 ( .A1(A[5]), .A2(B[5]), .ZN(n137) );
  XNOR2_X2 U164 ( .A(n143), .B(n17), .ZN(SUM[4]) );
  NAND2_X2 U168 ( .A1(n173), .A2(n142), .ZN(n17) );
  NAND2_X2 U171 ( .A1(A[4]), .A2(B[4]), .ZN(n142) );
  XNOR2_X2 U172 ( .A(n149), .B(n18), .ZN(SUM[3]) );
  NAND2_X2 U177 ( .A1(n174), .A2(n148), .ZN(n18) );
  NAND2_X2 U180 ( .A1(A[3]), .A2(B[3]), .ZN(n148) );
  XOR2_X2 U181 ( .A(n19), .B(n152), .Z(SUM[2]) );
  NAND2_X2 U183 ( .A1(n175), .A2(n151), .ZN(n19) );
  NAND2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n151) );
  XOR2_X2 U187 ( .A(n157), .B(n20), .Z(SUM[1]) );
  NAND2_X2 U190 ( .A1(n176), .A2(n155), .ZN(n20) );
  NAND2_X2 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n155) );
  NAND2_X2 U198 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  OR2_X2 U202 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  OR2_X4 U203 ( .A1(n30), .A2(n27), .ZN(n248) );
  AND2_X1 U204 ( .A1(n250), .A2(n157), .ZN(SUM[0]) );
  NOR2_X1 U205 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  OAI21_X1 U206 ( .B1(n114), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X1 U207 ( .B1(n86), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U208 ( .B1(n114), .B2(n56), .A(n57), .ZN(n55) );
  AOI21_X4 U209 ( .B1(n115), .B2(n47), .A(n48), .ZN(n1) );
  AOI21_X1 U210 ( .B1(n86), .B2(n67), .A(n68), .ZN(n66) );
  AOI21_X1 U211 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U212 ( .B1(n1), .B2(n37), .A(n38), .ZN(n36) );
  INV_X1 U213 ( .A(n40), .ZN(n38) );
  OAI21_X1 U214 ( .B1(n114), .B2(n101), .A(n102), .ZN(n100) );
  INV_X1 U215 ( .A(n104), .ZN(n102) );
  NOR2_X1 U216 ( .A1(n69), .A2(n60), .ZN(n58) );
  OAI21_X1 U217 ( .B1(n133), .B2(n125), .A(n128), .ZN(n124) );
  NOR2_X1 U218 ( .A1(n132), .A2(n125), .ZN(n123) );
  NOR2_X1 U219 ( .A1(n80), .A2(n73), .ZN(n67) );
  OAI21_X1 U220 ( .B1(n114), .B2(n94), .A(n95), .ZN(n93) );
  OAI21_X1 U221 ( .B1(n1), .B2(n44), .A(n45), .ZN(n43) );
  NOR2_X1 U222 ( .A1(n141), .A2(n136), .ZN(n130) );
  NOR2_X1 U223 ( .A1(n112), .A2(n109), .ZN(n103) );
  NOR2_X1 U224 ( .A1(n150), .A2(n147), .ZN(n145) );
  OAI21_X1 U225 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  OAI21_X1 U226 ( .B1(n120), .B2(n128), .A(n121), .ZN(n119) );
  NOR2_X1 U227 ( .A1(n44), .A2(n41), .ZN(n39) );
  NOR2_X1 U228 ( .A1(n98), .A2(n91), .ZN(n89) );
  NOR2_X1 U229 ( .A1(n60), .A2(n53), .ZN(n51) );
  OAI21_X1 U230 ( .B1(n31), .B2(n27), .A(n28), .ZN(n26) );
  NOR2_X1 U231 ( .A1(A[16]), .A2(B[16]), .ZN(n44) );
  NOR2_X1 U232 ( .A1(A[12]), .A2(B[12]), .ZN(n80) );
  NOR2_X1 U233 ( .A1(n83), .A2(n49), .ZN(n47) );
  OAI21_X2 U234 ( .B1(n84), .B2(n49), .A(n50), .ZN(n48) );
  OAI21_X1 U235 ( .B1(n1), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X1 U236 ( .B1(n114), .B2(n83), .A(n84), .ZN(n82) );
  OAI21_X1 U237 ( .B1(n114), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U238 ( .B1(n40), .B2(n247), .A(n33), .ZN(n31) );
  OAI21_X2 U239 ( .B1(n109), .B2(n113), .A(n110), .ZN(n104) );
  AOI21_X2 U240 ( .B1(n145), .B2(n153), .A(n146), .ZN(n144) );
  OAI21_X2 U241 ( .B1(n73), .B2(n81), .A(n74), .ZN(n68) );
  OAI21_X2 U242 ( .B1(n136), .B2(n142), .A(n137), .ZN(n131) );
  OAI21_X2 U243 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI21_X2 U244 ( .B1(n144), .B2(n116), .A(n117), .ZN(n115) );
  AOI21_X2 U245 ( .B1(n118), .B2(n131), .A(n119), .ZN(n117) );
  NOR2_X2 U246 ( .A1(n125), .A2(n120), .ZN(n118) );
  AOI21_X2 U247 ( .B1(n51), .B2(n68), .A(n52), .ZN(n50) );
  OAI21_X2 U248 ( .B1(n53), .B2(n63), .A(n54), .ZN(n52) );
  AOI21_X2 U249 ( .B1(n143), .B2(n123), .A(n124), .ZN(n122) );
  AOI21_X2 U250 ( .B1(n143), .B2(n173), .A(n140), .ZN(n138) );
  OAI21_X2 U251 ( .B1(n154), .B2(n157), .A(n155), .ZN(n153) );
  AOI21_X2 U252 ( .B1(n89), .B2(n104), .A(n90), .ZN(n84) );
  OAI21_X2 U253 ( .B1(n91), .B2(n99), .A(n92), .ZN(n90) );
  OAI21_X1 U254 ( .B1(n70), .B2(n60), .A(n63), .ZN(n59) );
  AOI21_X2 U255 ( .B1(n86), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X1 U256 ( .B1(n104), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U257 ( .B1(n114), .B2(n112), .A(n113), .ZN(n111) );
  OAI21_X1 U258 ( .B1(n152), .B2(n150), .A(n151), .ZN(n149) );
  NOR2_X2 U259 ( .A1(A[14]), .A2(B[14]), .ZN(n60) );
  NOR2_X2 U260 ( .A1(A[6]), .A2(B[6]), .ZN(n125) );
  NOR2_X2 U261 ( .A1(A[13]), .A2(B[13]), .ZN(n73) );
  NOR2_X2 U262 ( .A1(A[15]), .A2(B[15]), .ZN(n53) );
  NOR2_X2 U263 ( .A1(A[11]), .A2(B[11]), .ZN(n91) );
  NOR2_X2 U264 ( .A1(A[9]), .A2(B[9]), .ZN(n109) );
  NOR2_X2 U265 ( .A1(A[5]), .A2(B[5]), .ZN(n136) );
  NOR2_X2 U266 ( .A1(A[7]), .A2(B[7]), .ZN(n120) );
  NOR2_X2 U267 ( .A1(A[17]), .A2(B[17]), .ZN(n41) );
  NOR2_X2 U268 ( .A1(A[3]), .A2(B[3]), .ZN(n147) );
  NOR2_X2 U269 ( .A1(A[19]), .A2(B[19]), .ZN(n27) );
  NOR2_X1 U270 ( .A1(A[8]), .A2(B[8]), .ZN(n112) );
  NOR2_X2 U271 ( .A1(A[1]), .A2(B[1]), .ZN(n154) );
  NOR2_X1 U272 ( .A1(A[10]), .A2(B[10]), .ZN(n98) );
  NOR2_X1 U273 ( .A1(A[4]), .A2(B[4]), .ZN(n141) );
  OAI21_X2 U274 ( .B1(n1), .B2(n248), .A(n24), .ZN(SUM[20]) );
  OR2_X1 U275 ( .A1(A[0]), .A2(B[0]), .ZN(n250) );
  INV_X4 U276 ( .A(n99), .ZN(n97) );
  INV_X4 U277 ( .A(n84), .ZN(n86) );
  INV_X4 U278 ( .A(n83), .ZN(n85) );
  INV_X4 U279 ( .A(n81), .ZN(n79) );
  INV_X4 U280 ( .A(n68), .ZN(n70) );
  INV_X4 U281 ( .A(n67), .ZN(n69) );
  INV_X4 U282 ( .A(n39), .ZN(n37) );
  INV_X4 U283 ( .A(n35), .ZN(n33) );
  INV_X4 U284 ( .A(n26), .ZN(n24) );
  INV_X4 U285 ( .A(n154), .ZN(n176) );
  INV_X4 U286 ( .A(n150), .ZN(n175) );
  INV_X4 U287 ( .A(n147), .ZN(n174) );
  INV_X4 U288 ( .A(n136), .ZN(n172) );
  INV_X4 U289 ( .A(n125), .ZN(n171) );
  INV_X4 U290 ( .A(n120), .ZN(n170) );
  INV_X4 U291 ( .A(n112), .ZN(n169) );
  INV_X4 U292 ( .A(n109), .ZN(n168) );
  INV_X4 U293 ( .A(n98), .ZN(n96) );
  INV_X4 U294 ( .A(n91), .ZN(n166) );
  INV_X4 U295 ( .A(n80), .ZN(n78) );
  INV_X4 U296 ( .A(n73), .ZN(n164) );
  INV_X4 U297 ( .A(n60), .ZN(n163) );
  INV_X4 U298 ( .A(n53), .ZN(n162) );
  INV_X4 U299 ( .A(n44), .ZN(n161) );
  INV_X4 U300 ( .A(n41), .ZN(n160) );
  INV_X4 U301 ( .A(n27), .ZN(n158) );
  INV_X4 U302 ( .A(n153), .ZN(n152) );
  INV_X4 U303 ( .A(n144), .ZN(n143) );
  INV_X4 U304 ( .A(n142), .ZN(n140) );
  INV_X4 U305 ( .A(n141), .ZN(n173) );
  INV_X4 U306 ( .A(n131), .ZN(n133) );
  INV_X4 U307 ( .A(n130), .ZN(n132) );
  INV_X4 U308 ( .A(n115), .ZN(n114) );
  INV_X4 U309 ( .A(n103), .ZN(n101) );
endmodule


module pipleline_stage_6 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n106;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;

  pipleline_stage_6_DW01_add_1 add_268 ( .A({1'b0, divided[26:7]}), .B({1'b0, 
        divisor}), .CI(1'b0), .SUM(stage_result) );
  BUF_X4 U5 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U6 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U7 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U8 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U9 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U10 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U11 ( .A(divided[0]), .Z(stage_out[1]) );
  INV_X16 U12 ( .A(n106), .ZN(q) );
  XNOR2_X2 U13 ( .A(divided[27]), .B(stage_result[20]), .ZN(n106) );
  MUX2_X2 U14 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U15 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U16 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U17 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U18 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U19 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U20 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U21 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U22 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U23 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U24 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U25 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U26 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U27 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U28 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U29 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U30 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U31 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U32 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U33 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64, n65,
         n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n128, n129, n130, n131, n132, n133, n136, n137, n138, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n157, n158, n160, n161, n162, n163, n164,
         n166, n168, n169, n170, n171, n172, n173, n174, n175, n176, n247,
         n249;

  XNOR2_X2 U3 ( .A(n29), .B(n2), .ZN(SUM[19]) );
  NAND2_X2 U9 ( .A1(n158), .A2(n28), .ZN(n2) );
  NAND2_X2 U12 ( .A1(A[19]), .A2(B[19]), .ZN(n28) );
  XNOR2_X2 U13 ( .A(n36), .B(n3), .ZN(SUM[18]) );
  NAND2_X2 U15 ( .A1(n39), .A2(n32), .ZN(n30) );
  NAND2_X2 U19 ( .A1(n32), .A2(n35), .ZN(n3) );
  NAND2_X2 U22 ( .A1(A[18]), .A2(B[18]), .ZN(n35) );
  XNOR2_X2 U23 ( .A(n43), .B(n4), .ZN(SUM[17]) );
  NAND2_X2 U29 ( .A1(n160), .A2(n42), .ZN(n4) );
  NAND2_X2 U32 ( .A1(A[17]), .A2(B[17]), .ZN(n42) );
  XOR2_X2 U33 ( .A(n5), .B(n1), .Z(SUM[16]) );
  NAND2_X2 U35 ( .A1(n161), .A2(n45), .ZN(n5) );
  NAND2_X2 U38 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U39 ( .A(n55), .B(n6), .ZN(SUM[15]) );
  NAND2_X2 U43 ( .A1(n67), .A2(n51), .ZN(n49) );
  NAND2_X2 U47 ( .A1(n162), .A2(n54), .ZN(n6) );
  NAND2_X2 U50 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  XNOR2_X2 U51 ( .A(n64), .B(n7), .ZN(SUM[14]) );
  NAND2_X2 U53 ( .A1(n58), .A2(n85), .ZN(n56) );
  NAND2_X2 U59 ( .A1(n163), .A2(n63), .ZN(n7) );
  NAND2_X2 U62 ( .A1(A[14]), .A2(B[14]), .ZN(n63) );
  XNOR2_X2 U63 ( .A(n75), .B(n8), .ZN(SUM[13]) );
  NAND2_X2 U65 ( .A1(n85), .A2(n67), .ZN(n65) );
  NAND2_X2 U73 ( .A1(n164), .A2(n74), .ZN(n8) );
  NAND2_X2 U76 ( .A1(A[13]), .A2(B[13]), .ZN(n74) );
  XNOR2_X2 U77 ( .A(n82), .B(n9), .ZN(SUM[12]) );
  NAND2_X2 U79 ( .A1(n85), .A2(n78), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n78), .A2(n81), .ZN(n9) );
  NAND2_X2 U86 ( .A1(A[12]), .A2(B[12]), .ZN(n81) );
  XNOR2_X2 U87 ( .A(n93), .B(n10), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(n103), .A2(n89), .ZN(n83) );
  NAND2_X2 U97 ( .A1(n166), .A2(n92), .ZN(n10) );
  NAND2_X2 U100 ( .A1(A[11]), .A2(B[11]), .ZN(n92) );
  XNOR2_X2 U101 ( .A(n100), .B(n11), .ZN(SUM[10]) );
  NAND2_X2 U103 ( .A1(n103), .A2(n96), .ZN(n94) );
  NAND2_X2 U107 ( .A1(n96), .A2(n99), .ZN(n11) );
  NAND2_X2 U110 ( .A1(A[10]), .A2(B[10]), .ZN(n99) );
  XNOR2_X2 U111 ( .A(n111), .B(n12), .ZN(SUM[9]) );
  NAND2_X2 U121 ( .A1(n168), .A2(n110), .ZN(n12) );
  NAND2_X2 U124 ( .A1(A[9]), .A2(B[9]), .ZN(n110) );
  XOR2_X2 U125 ( .A(n13), .B(n114), .Z(SUM[8]) );
  NAND2_X2 U127 ( .A1(n169), .A2(n113), .ZN(n13) );
  NAND2_X2 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n113) );
  XOR2_X2 U131 ( .A(n14), .B(n122), .Z(SUM[7]) );
  NAND2_X2 U134 ( .A1(n130), .A2(n118), .ZN(n116) );
  NAND2_X2 U138 ( .A1(n170), .A2(n121), .ZN(n14) );
  NAND2_X2 U141 ( .A1(A[7]), .A2(B[7]), .ZN(n121) );
  XOR2_X2 U142 ( .A(n15), .B(n129), .Z(SUM[6]) );
  NAND2_X2 U148 ( .A1(n171), .A2(n128), .ZN(n15) );
  NAND2_X2 U151 ( .A1(A[6]), .A2(B[6]), .ZN(n128) );
  XOR2_X2 U152 ( .A(n16), .B(n138), .Z(SUM[5]) );
  NAND2_X2 U160 ( .A1(n172), .A2(n137), .ZN(n16) );
  NAND2_X2 U163 ( .A1(A[5]), .A2(B[5]), .ZN(n137) );
  XNOR2_X2 U164 ( .A(n143), .B(n17), .ZN(SUM[4]) );
  NAND2_X2 U168 ( .A1(n173), .A2(n142), .ZN(n17) );
  NAND2_X2 U171 ( .A1(A[4]), .A2(B[4]), .ZN(n142) );
  XNOR2_X2 U172 ( .A(n149), .B(n18), .ZN(SUM[3]) );
  NAND2_X2 U177 ( .A1(n174), .A2(n148), .ZN(n18) );
  NAND2_X2 U180 ( .A1(A[3]), .A2(B[3]), .ZN(n148) );
  XOR2_X2 U181 ( .A(n19), .B(n152), .Z(SUM[2]) );
  NAND2_X2 U183 ( .A1(n175), .A2(n151), .ZN(n19) );
  NAND2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n151) );
  XOR2_X2 U187 ( .A(n157), .B(n20), .Z(SUM[1]) );
  NAND2_X2 U190 ( .A1(n176), .A2(n155), .ZN(n20) );
  NAND2_X2 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n155) );
  NAND2_X2 U198 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  OR2_X4 U202 ( .A1(n30), .A2(n27), .ZN(n247) );
  AND2_X1 U203 ( .A1(n249), .A2(n157), .ZN(SUM[0]) );
  NOR2_X1 U204 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  NOR2_X1 U205 ( .A1(A[18]), .A2(B[18]), .ZN(n34) );
  OAI21_X1 U206 ( .B1(n114), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X1 U207 ( .B1(n86), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U208 ( .B1(n114), .B2(n56), .A(n57), .ZN(n55) );
  AOI21_X4 U209 ( .B1(n115), .B2(n47), .A(n48), .ZN(n1) );
  AOI21_X1 U210 ( .B1(n86), .B2(n67), .A(n68), .ZN(n66) );
  AOI21_X1 U211 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U212 ( .B1(n1), .B2(n37), .A(n38), .ZN(n36) );
  INV_X1 U213 ( .A(n40), .ZN(n38) );
  OAI21_X1 U214 ( .B1(n114), .B2(n101), .A(n102), .ZN(n100) );
  INV_X1 U215 ( .A(n104), .ZN(n102) );
  NOR2_X1 U216 ( .A1(n69), .A2(n60), .ZN(n58) );
  OAI21_X1 U217 ( .B1(n133), .B2(n125), .A(n128), .ZN(n124) );
  NOR2_X1 U218 ( .A1(n132), .A2(n125), .ZN(n123) );
  NOR2_X1 U219 ( .A1(n80), .A2(n73), .ZN(n67) );
  OAI21_X1 U220 ( .B1(n114), .B2(n94), .A(n95), .ZN(n93) );
  OAI21_X1 U221 ( .B1(n1), .B2(n44), .A(n45), .ZN(n43) );
  NOR2_X1 U222 ( .A1(n141), .A2(n136), .ZN(n130) );
  NOR2_X1 U223 ( .A1(n112), .A2(n109), .ZN(n103) );
  NOR2_X1 U224 ( .A1(n150), .A2(n147), .ZN(n145) );
  OAI21_X1 U225 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  OAI21_X1 U226 ( .B1(n120), .B2(n128), .A(n121), .ZN(n119) );
  NOR2_X1 U227 ( .A1(n44), .A2(n41), .ZN(n39) );
  NOR2_X1 U228 ( .A1(n98), .A2(n91), .ZN(n89) );
  NOR2_X1 U229 ( .A1(n60), .A2(n53), .ZN(n51) );
  OAI21_X1 U230 ( .B1(n31), .B2(n27), .A(n28), .ZN(n26) );
  NOR2_X1 U231 ( .A1(A[16]), .A2(B[16]), .ZN(n44) );
  NOR2_X1 U232 ( .A1(A[12]), .A2(B[12]), .ZN(n80) );
  NOR2_X1 U233 ( .A1(n83), .A2(n49), .ZN(n47) );
  OAI21_X2 U234 ( .B1(n84), .B2(n49), .A(n50), .ZN(n48) );
  OAI21_X1 U235 ( .B1(n1), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X1 U236 ( .B1(n114), .B2(n83), .A(n84), .ZN(n82) );
  OAI21_X1 U237 ( .B1(n114), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U238 ( .B1(n40), .B2(n32), .A(n33), .ZN(n31) );
  OAI21_X2 U239 ( .B1(n109), .B2(n113), .A(n110), .ZN(n104) );
  AOI21_X2 U240 ( .B1(n145), .B2(n153), .A(n146), .ZN(n144) );
  OAI21_X2 U241 ( .B1(n73), .B2(n81), .A(n74), .ZN(n68) );
  OAI21_X2 U242 ( .B1(n136), .B2(n142), .A(n137), .ZN(n131) );
  OAI21_X2 U243 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI21_X2 U244 ( .B1(n144), .B2(n116), .A(n117), .ZN(n115) );
  AOI21_X2 U245 ( .B1(n118), .B2(n131), .A(n119), .ZN(n117) );
  NOR2_X2 U246 ( .A1(n125), .A2(n120), .ZN(n118) );
  AOI21_X2 U247 ( .B1(n51), .B2(n68), .A(n52), .ZN(n50) );
  OAI21_X2 U248 ( .B1(n53), .B2(n63), .A(n54), .ZN(n52) );
  AOI21_X2 U249 ( .B1(n143), .B2(n123), .A(n124), .ZN(n122) );
  AOI21_X2 U250 ( .B1(n143), .B2(n173), .A(n140), .ZN(n138) );
  OAI21_X2 U251 ( .B1(n154), .B2(n157), .A(n155), .ZN(n153) );
  AOI21_X2 U252 ( .B1(n89), .B2(n104), .A(n90), .ZN(n84) );
  OAI21_X2 U253 ( .B1(n91), .B2(n99), .A(n92), .ZN(n90) );
  OAI21_X1 U254 ( .B1(n70), .B2(n60), .A(n63), .ZN(n59) );
  AOI21_X2 U255 ( .B1(n86), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X1 U256 ( .B1(n104), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U257 ( .B1(n114), .B2(n112), .A(n113), .ZN(n111) );
  OAI21_X1 U258 ( .B1(n152), .B2(n150), .A(n151), .ZN(n149) );
  NOR2_X2 U259 ( .A1(A[14]), .A2(B[14]), .ZN(n60) );
  NOR2_X2 U260 ( .A1(A[6]), .A2(B[6]), .ZN(n125) );
  NOR2_X2 U261 ( .A1(A[13]), .A2(B[13]), .ZN(n73) );
  NOR2_X2 U262 ( .A1(A[15]), .A2(B[15]), .ZN(n53) );
  NOR2_X2 U263 ( .A1(A[11]), .A2(B[11]), .ZN(n91) );
  NOR2_X2 U264 ( .A1(A[9]), .A2(B[9]), .ZN(n109) );
  NOR2_X2 U265 ( .A1(A[5]), .A2(B[5]), .ZN(n136) );
  NOR2_X2 U266 ( .A1(A[7]), .A2(B[7]), .ZN(n120) );
  NOR2_X2 U267 ( .A1(A[17]), .A2(B[17]), .ZN(n41) );
  NOR2_X2 U268 ( .A1(A[3]), .A2(B[3]), .ZN(n147) );
  NOR2_X2 U269 ( .A1(A[19]), .A2(B[19]), .ZN(n27) );
  NOR2_X1 U270 ( .A1(A[8]), .A2(B[8]), .ZN(n112) );
  NOR2_X2 U271 ( .A1(A[1]), .A2(B[1]), .ZN(n154) );
  NOR2_X1 U272 ( .A1(A[10]), .A2(B[10]), .ZN(n98) );
  NOR2_X1 U273 ( .A1(A[4]), .A2(B[4]), .ZN(n141) );
  OAI21_X2 U274 ( .B1(n1), .B2(n247), .A(n24), .ZN(SUM[20]) );
  OR2_X1 U275 ( .A1(A[0]), .A2(B[0]), .ZN(n249) );
  INV_X4 U276 ( .A(n99), .ZN(n97) );
  INV_X4 U277 ( .A(n84), .ZN(n86) );
  INV_X4 U278 ( .A(n83), .ZN(n85) );
  INV_X4 U279 ( .A(n81), .ZN(n79) );
  INV_X4 U280 ( .A(n68), .ZN(n70) );
  INV_X4 U281 ( .A(n67), .ZN(n69) );
  INV_X4 U282 ( .A(n39), .ZN(n37) );
  INV_X4 U283 ( .A(n35), .ZN(n33) );
  INV_X4 U284 ( .A(n26), .ZN(n24) );
  INV_X4 U285 ( .A(n154), .ZN(n176) );
  INV_X4 U286 ( .A(n150), .ZN(n175) );
  INV_X4 U287 ( .A(n147), .ZN(n174) );
  INV_X4 U288 ( .A(n136), .ZN(n172) );
  INV_X4 U289 ( .A(n125), .ZN(n171) );
  INV_X4 U290 ( .A(n120), .ZN(n170) );
  INV_X4 U291 ( .A(n112), .ZN(n169) );
  INV_X4 U292 ( .A(n109), .ZN(n168) );
  INV_X4 U293 ( .A(n98), .ZN(n96) );
  INV_X4 U294 ( .A(n91), .ZN(n166) );
  INV_X4 U295 ( .A(n80), .ZN(n78) );
  INV_X4 U296 ( .A(n73), .ZN(n164) );
  INV_X4 U297 ( .A(n60), .ZN(n163) );
  INV_X4 U298 ( .A(n53), .ZN(n162) );
  INV_X4 U299 ( .A(n44), .ZN(n161) );
  INV_X4 U300 ( .A(n41), .ZN(n160) );
  INV_X4 U301 ( .A(n34), .ZN(n32) );
  INV_X4 U302 ( .A(n27), .ZN(n158) );
  INV_X4 U303 ( .A(n153), .ZN(n152) );
  INV_X4 U304 ( .A(n144), .ZN(n143) );
  INV_X4 U305 ( .A(n142), .ZN(n140) );
  INV_X4 U306 ( .A(n141), .ZN(n173) );
  INV_X4 U307 ( .A(n131), .ZN(n133) );
  INV_X4 U308 ( .A(n130), .ZN(n132) );
  INV_X4 U309 ( .A(n115), .ZN(n114) );
  INV_X4 U310 ( .A(n103), .ZN(n101) );
endmodule


module pipleline_stage_5 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n106;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;

  pipleline_stage_5_DW01_add_1 add_268 ( .A({1'b0, divided[26:7]}), .B({1'b0, 
        divisor}), .CI(1'b0), .SUM(stage_result) );
  BUF_X4 U5 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U6 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U7 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U8 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U9 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U10 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U11 ( .A(divided[0]), .Z(stage_out[1]) );
  INV_X16 U12 ( .A(n106), .ZN(q) );
  XNOR2_X2 U13 ( .A(divided[27]), .B(stage_result[20]), .ZN(n106) );
  MUX2_X2 U14 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U15 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U16 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U17 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U18 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U19 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U20 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U21 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U22 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U23 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U24 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U25 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U26 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U27 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U28 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U29 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U30 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U31 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U32 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U33 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n24, n26, n27, n28, n29, n30, n31, n33, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64, n65, n66, n67,
         n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n128, n129, n130, n131, n132, n133, n136, n137, n138, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n157, n158, n160, n161, n162, n163, n164, n166,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n247, n248,
         n250;

  XNOR2_X2 U3 ( .A(n29), .B(n2), .ZN(SUM[19]) );
  NAND2_X2 U9 ( .A1(n158), .A2(n28), .ZN(n2) );
  NAND2_X2 U12 ( .A1(A[19]), .A2(B[19]), .ZN(n28) );
  XNOR2_X2 U13 ( .A(n36), .B(n3), .ZN(SUM[18]) );
  NAND2_X2 U15 ( .A1(n39), .A2(n247), .ZN(n30) );
  NAND2_X2 U19 ( .A1(n247), .A2(n35), .ZN(n3) );
  NAND2_X2 U22 ( .A1(A[18]), .A2(B[18]), .ZN(n35) );
  XNOR2_X2 U23 ( .A(n43), .B(n4), .ZN(SUM[17]) );
  NAND2_X2 U29 ( .A1(n160), .A2(n42), .ZN(n4) );
  NAND2_X2 U32 ( .A1(A[17]), .A2(B[17]), .ZN(n42) );
  XOR2_X2 U33 ( .A(n5), .B(n1), .Z(SUM[16]) );
  NAND2_X2 U35 ( .A1(n161), .A2(n45), .ZN(n5) );
  NAND2_X2 U38 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U39 ( .A(n55), .B(n6), .ZN(SUM[15]) );
  NAND2_X2 U43 ( .A1(n67), .A2(n51), .ZN(n49) );
  NAND2_X2 U47 ( .A1(n162), .A2(n54), .ZN(n6) );
  NAND2_X2 U50 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  XNOR2_X2 U51 ( .A(n64), .B(n7), .ZN(SUM[14]) );
  NAND2_X2 U53 ( .A1(n58), .A2(n85), .ZN(n56) );
  NAND2_X2 U59 ( .A1(n163), .A2(n63), .ZN(n7) );
  NAND2_X2 U62 ( .A1(A[14]), .A2(B[14]), .ZN(n63) );
  XNOR2_X2 U63 ( .A(n75), .B(n8), .ZN(SUM[13]) );
  NAND2_X2 U65 ( .A1(n85), .A2(n67), .ZN(n65) );
  NAND2_X2 U73 ( .A1(n164), .A2(n74), .ZN(n8) );
  NAND2_X2 U76 ( .A1(A[13]), .A2(B[13]), .ZN(n74) );
  XNOR2_X2 U77 ( .A(n82), .B(n9), .ZN(SUM[12]) );
  NAND2_X2 U79 ( .A1(n85), .A2(n78), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n78), .A2(n81), .ZN(n9) );
  NAND2_X2 U86 ( .A1(A[12]), .A2(B[12]), .ZN(n81) );
  XNOR2_X2 U87 ( .A(n93), .B(n10), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(n103), .A2(n89), .ZN(n83) );
  NAND2_X2 U97 ( .A1(n166), .A2(n92), .ZN(n10) );
  NAND2_X2 U100 ( .A1(A[11]), .A2(B[11]), .ZN(n92) );
  XNOR2_X2 U101 ( .A(n100), .B(n11), .ZN(SUM[10]) );
  NAND2_X2 U103 ( .A1(n103), .A2(n96), .ZN(n94) );
  NAND2_X2 U107 ( .A1(n96), .A2(n99), .ZN(n11) );
  NAND2_X2 U110 ( .A1(A[10]), .A2(B[10]), .ZN(n99) );
  XNOR2_X2 U111 ( .A(n111), .B(n12), .ZN(SUM[9]) );
  NAND2_X2 U121 ( .A1(n168), .A2(n110), .ZN(n12) );
  NAND2_X2 U124 ( .A1(A[9]), .A2(B[9]), .ZN(n110) );
  XOR2_X2 U125 ( .A(n13), .B(n114), .Z(SUM[8]) );
  NAND2_X2 U127 ( .A1(n169), .A2(n113), .ZN(n13) );
  NAND2_X2 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n113) );
  XOR2_X2 U131 ( .A(n14), .B(n122), .Z(SUM[7]) );
  NAND2_X2 U134 ( .A1(n130), .A2(n118), .ZN(n116) );
  NAND2_X2 U138 ( .A1(n170), .A2(n121), .ZN(n14) );
  NAND2_X2 U141 ( .A1(A[7]), .A2(B[7]), .ZN(n121) );
  XOR2_X2 U142 ( .A(n15), .B(n129), .Z(SUM[6]) );
  NAND2_X2 U148 ( .A1(n171), .A2(n128), .ZN(n15) );
  NAND2_X2 U151 ( .A1(A[6]), .A2(B[6]), .ZN(n128) );
  XOR2_X2 U152 ( .A(n16), .B(n138), .Z(SUM[5]) );
  NAND2_X2 U160 ( .A1(n172), .A2(n137), .ZN(n16) );
  NAND2_X2 U163 ( .A1(A[5]), .A2(B[5]), .ZN(n137) );
  XNOR2_X2 U164 ( .A(n143), .B(n17), .ZN(SUM[4]) );
  NAND2_X2 U168 ( .A1(n173), .A2(n142), .ZN(n17) );
  NAND2_X2 U171 ( .A1(A[4]), .A2(B[4]), .ZN(n142) );
  XNOR2_X2 U172 ( .A(n149), .B(n18), .ZN(SUM[3]) );
  NAND2_X2 U177 ( .A1(n174), .A2(n148), .ZN(n18) );
  NAND2_X2 U180 ( .A1(A[3]), .A2(B[3]), .ZN(n148) );
  XOR2_X2 U181 ( .A(n19), .B(n152), .Z(SUM[2]) );
  NAND2_X2 U183 ( .A1(n175), .A2(n151), .ZN(n19) );
  NAND2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n151) );
  XOR2_X2 U187 ( .A(n157), .B(n20), .Z(SUM[1]) );
  NAND2_X2 U190 ( .A1(n176), .A2(n155), .ZN(n20) );
  NAND2_X2 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n155) );
  NAND2_X2 U198 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  OR2_X2 U202 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  OR2_X4 U203 ( .A1(n30), .A2(n27), .ZN(n248) );
  AND2_X1 U204 ( .A1(n250), .A2(n157), .ZN(SUM[0]) );
  NOR2_X1 U205 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  OAI21_X1 U206 ( .B1(n114), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X1 U207 ( .B1(n86), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U208 ( .B1(n114), .B2(n56), .A(n57), .ZN(n55) );
  AOI21_X4 U209 ( .B1(n115), .B2(n47), .A(n48), .ZN(n1) );
  AOI21_X1 U210 ( .B1(n86), .B2(n67), .A(n68), .ZN(n66) );
  AOI21_X1 U211 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U212 ( .B1(n1), .B2(n37), .A(n38), .ZN(n36) );
  INV_X1 U213 ( .A(n40), .ZN(n38) );
  OAI21_X1 U214 ( .B1(n114), .B2(n101), .A(n102), .ZN(n100) );
  INV_X1 U215 ( .A(n104), .ZN(n102) );
  NOR2_X1 U216 ( .A1(n69), .A2(n60), .ZN(n58) );
  OAI21_X1 U217 ( .B1(n133), .B2(n125), .A(n128), .ZN(n124) );
  NOR2_X1 U218 ( .A1(n132), .A2(n125), .ZN(n123) );
  NOR2_X1 U219 ( .A1(n80), .A2(n73), .ZN(n67) );
  OAI21_X1 U220 ( .B1(n114), .B2(n94), .A(n95), .ZN(n93) );
  OAI21_X1 U221 ( .B1(n1), .B2(n44), .A(n45), .ZN(n43) );
  NOR2_X1 U222 ( .A1(n141), .A2(n136), .ZN(n130) );
  NOR2_X1 U223 ( .A1(n112), .A2(n109), .ZN(n103) );
  NOR2_X1 U224 ( .A1(n150), .A2(n147), .ZN(n145) );
  OAI21_X1 U225 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  OAI21_X1 U226 ( .B1(n120), .B2(n128), .A(n121), .ZN(n119) );
  NOR2_X1 U227 ( .A1(n44), .A2(n41), .ZN(n39) );
  NOR2_X1 U228 ( .A1(n98), .A2(n91), .ZN(n89) );
  NOR2_X1 U229 ( .A1(n60), .A2(n53), .ZN(n51) );
  OAI21_X1 U230 ( .B1(n31), .B2(n27), .A(n28), .ZN(n26) );
  NOR2_X1 U231 ( .A1(A[16]), .A2(B[16]), .ZN(n44) );
  NOR2_X1 U232 ( .A1(A[12]), .A2(B[12]), .ZN(n80) );
  NOR2_X1 U233 ( .A1(n83), .A2(n49), .ZN(n47) );
  OAI21_X2 U234 ( .B1(n84), .B2(n49), .A(n50), .ZN(n48) );
  OAI21_X1 U235 ( .B1(n1), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X1 U236 ( .B1(n114), .B2(n83), .A(n84), .ZN(n82) );
  OAI21_X1 U237 ( .B1(n114), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U238 ( .B1(n40), .B2(n247), .A(n33), .ZN(n31) );
  OAI21_X2 U239 ( .B1(n109), .B2(n113), .A(n110), .ZN(n104) );
  AOI21_X2 U240 ( .B1(n145), .B2(n153), .A(n146), .ZN(n144) );
  OAI21_X2 U241 ( .B1(n73), .B2(n81), .A(n74), .ZN(n68) );
  OAI21_X2 U242 ( .B1(n136), .B2(n142), .A(n137), .ZN(n131) );
  OAI21_X2 U243 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI21_X2 U244 ( .B1(n144), .B2(n116), .A(n117), .ZN(n115) );
  AOI21_X2 U245 ( .B1(n118), .B2(n131), .A(n119), .ZN(n117) );
  NOR2_X2 U246 ( .A1(n125), .A2(n120), .ZN(n118) );
  AOI21_X2 U247 ( .B1(n51), .B2(n68), .A(n52), .ZN(n50) );
  OAI21_X2 U248 ( .B1(n53), .B2(n63), .A(n54), .ZN(n52) );
  AOI21_X2 U249 ( .B1(n143), .B2(n123), .A(n124), .ZN(n122) );
  AOI21_X2 U250 ( .B1(n143), .B2(n173), .A(n140), .ZN(n138) );
  OAI21_X2 U251 ( .B1(n154), .B2(n157), .A(n155), .ZN(n153) );
  AOI21_X2 U252 ( .B1(n89), .B2(n104), .A(n90), .ZN(n84) );
  OAI21_X2 U253 ( .B1(n91), .B2(n99), .A(n92), .ZN(n90) );
  OAI21_X1 U254 ( .B1(n70), .B2(n60), .A(n63), .ZN(n59) );
  AOI21_X2 U255 ( .B1(n86), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X1 U256 ( .B1(n104), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U257 ( .B1(n114), .B2(n112), .A(n113), .ZN(n111) );
  OAI21_X1 U258 ( .B1(n152), .B2(n150), .A(n151), .ZN(n149) );
  NOR2_X2 U259 ( .A1(A[14]), .A2(B[14]), .ZN(n60) );
  NOR2_X2 U260 ( .A1(A[6]), .A2(B[6]), .ZN(n125) );
  NOR2_X2 U261 ( .A1(A[13]), .A2(B[13]), .ZN(n73) );
  NOR2_X2 U262 ( .A1(A[15]), .A2(B[15]), .ZN(n53) );
  NOR2_X2 U263 ( .A1(A[11]), .A2(B[11]), .ZN(n91) );
  NOR2_X2 U264 ( .A1(A[9]), .A2(B[9]), .ZN(n109) );
  NOR2_X2 U265 ( .A1(A[5]), .A2(B[5]), .ZN(n136) );
  NOR2_X2 U266 ( .A1(A[7]), .A2(B[7]), .ZN(n120) );
  NOR2_X2 U267 ( .A1(A[17]), .A2(B[17]), .ZN(n41) );
  NOR2_X2 U268 ( .A1(A[3]), .A2(B[3]), .ZN(n147) );
  NOR2_X2 U269 ( .A1(A[19]), .A2(B[19]), .ZN(n27) );
  NOR2_X1 U270 ( .A1(A[8]), .A2(B[8]), .ZN(n112) );
  NOR2_X2 U271 ( .A1(A[1]), .A2(B[1]), .ZN(n154) );
  NOR2_X1 U272 ( .A1(A[10]), .A2(B[10]), .ZN(n98) );
  NOR2_X1 U273 ( .A1(A[4]), .A2(B[4]), .ZN(n141) );
  OAI21_X2 U274 ( .B1(n1), .B2(n248), .A(n24), .ZN(SUM[20]) );
  OR2_X1 U275 ( .A1(A[0]), .A2(B[0]), .ZN(n250) );
  INV_X4 U276 ( .A(n99), .ZN(n97) );
  INV_X4 U277 ( .A(n84), .ZN(n86) );
  INV_X4 U278 ( .A(n83), .ZN(n85) );
  INV_X4 U279 ( .A(n81), .ZN(n79) );
  INV_X4 U280 ( .A(n68), .ZN(n70) );
  INV_X4 U281 ( .A(n67), .ZN(n69) );
  INV_X4 U282 ( .A(n39), .ZN(n37) );
  INV_X4 U283 ( .A(n35), .ZN(n33) );
  INV_X4 U284 ( .A(n26), .ZN(n24) );
  INV_X4 U285 ( .A(n154), .ZN(n176) );
  INV_X4 U286 ( .A(n150), .ZN(n175) );
  INV_X4 U287 ( .A(n147), .ZN(n174) );
  INV_X4 U288 ( .A(n136), .ZN(n172) );
  INV_X4 U289 ( .A(n125), .ZN(n171) );
  INV_X4 U290 ( .A(n120), .ZN(n170) );
  INV_X4 U291 ( .A(n112), .ZN(n169) );
  INV_X4 U292 ( .A(n109), .ZN(n168) );
  INV_X4 U293 ( .A(n98), .ZN(n96) );
  INV_X4 U294 ( .A(n91), .ZN(n166) );
  INV_X4 U295 ( .A(n80), .ZN(n78) );
  INV_X4 U296 ( .A(n73), .ZN(n164) );
  INV_X4 U297 ( .A(n60), .ZN(n163) );
  INV_X4 U298 ( .A(n53), .ZN(n162) );
  INV_X4 U299 ( .A(n44), .ZN(n161) );
  INV_X4 U300 ( .A(n41), .ZN(n160) );
  INV_X4 U301 ( .A(n27), .ZN(n158) );
  INV_X4 U302 ( .A(n153), .ZN(n152) );
  INV_X4 U303 ( .A(n144), .ZN(n143) );
  INV_X4 U304 ( .A(n142), .ZN(n140) );
  INV_X4 U305 ( .A(n141), .ZN(n173) );
  INV_X4 U306 ( .A(n131), .ZN(n133) );
  INV_X4 U307 ( .A(n130), .ZN(n132) );
  INV_X4 U308 ( .A(n115), .ZN(n114) );
  INV_X4 U309 ( .A(n103), .ZN(n101) );
endmodule


module pipleline_stage_4 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n106;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;

  pipleline_stage_4_DW01_add_1 add_268 ( .A({1'b0, divided[26:7]}), .B({1'b0, 
        divisor}), .CI(1'b0), .SUM(stage_result) );
  BUF_X4 U5 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U6 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U7 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U8 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U9 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U10 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U11 ( .A(divided[0]), .Z(stage_out[1]) );
  INV_X16 U12 ( .A(n106), .ZN(q) );
  XNOR2_X2 U13 ( .A(divided[27]), .B(stage_result[20]), .ZN(n106) );
  MUX2_X2 U14 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U15 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U16 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U17 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U18 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U19 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U20 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U21 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U22 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U23 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U24 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U25 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U26 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U27 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U28 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U29 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U30 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U31 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U32 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U33 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64, n65,
         n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n128, n129, n130, n131, n132, n133, n136, n137, n138, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n157, n158, n160, n161, n162, n163, n164,
         n166, n168, n169, n170, n171, n172, n173, n174, n175, n176, n247,
         n249;

  XNOR2_X2 U3 ( .A(n29), .B(n2), .ZN(SUM[19]) );
  NAND2_X2 U9 ( .A1(n158), .A2(n28), .ZN(n2) );
  NAND2_X2 U12 ( .A1(A[19]), .A2(B[19]), .ZN(n28) );
  XNOR2_X2 U13 ( .A(n36), .B(n3), .ZN(SUM[18]) );
  NAND2_X2 U15 ( .A1(n39), .A2(n32), .ZN(n30) );
  NAND2_X2 U19 ( .A1(n32), .A2(n35), .ZN(n3) );
  NAND2_X2 U22 ( .A1(A[18]), .A2(B[18]), .ZN(n35) );
  XNOR2_X2 U23 ( .A(n43), .B(n4), .ZN(SUM[17]) );
  NAND2_X2 U29 ( .A1(n160), .A2(n42), .ZN(n4) );
  NAND2_X2 U32 ( .A1(A[17]), .A2(B[17]), .ZN(n42) );
  XOR2_X2 U33 ( .A(n5), .B(n1), .Z(SUM[16]) );
  NAND2_X2 U35 ( .A1(n161), .A2(n45), .ZN(n5) );
  NAND2_X2 U38 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U39 ( .A(n55), .B(n6), .ZN(SUM[15]) );
  NAND2_X2 U43 ( .A1(n67), .A2(n51), .ZN(n49) );
  NAND2_X2 U47 ( .A1(n162), .A2(n54), .ZN(n6) );
  NAND2_X2 U50 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  XNOR2_X2 U51 ( .A(n64), .B(n7), .ZN(SUM[14]) );
  NAND2_X2 U53 ( .A1(n58), .A2(n85), .ZN(n56) );
  NAND2_X2 U59 ( .A1(n163), .A2(n63), .ZN(n7) );
  NAND2_X2 U62 ( .A1(A[14]), .A2(B[14]), .ZN(n63) );
  XNOR2_X2 U63 ( .A(n75), .B(n8), .ZN(SUM[13]) );
  NAND2_X2 U65 ( .A1(n85), .A2(n67), .ZN(n65) );
  NAND2_X2 U73 ( .A1(n164), .A2(n74), .ZN(n8) );
  NAND2_X2 U76 ( .A1(A[13]), .A2(B[13]), .ZN(n74) );
  XNOR2_X2 U77 ( .A(n82), .B(n9), .ZN(SUM[12]) );
  NAND2_X2 U79 ( .A1(n85), .A2(n78), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n78), .A2(n81), .ZN(n9) );
  NAND2_X2 U86 ( .A1(A[12]), .A2(B[12]), .ZN(n81) );
  XNOR2_X2 U87 ( .A(n93), .B(n10), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(n103), .A2(n89), .ZN(n83) );
  NAND2_X2 U97 ( .A1(n166), .A2(n92), .ZN(n10) );
  NAND2_X2 U100 ( .A1(A[11]), .A2(B[11]), .ZN(n92) );
  XNOR2_X2 U101 ( .A(n100), .B(n11), .ZN(SUM[10]) );
  NAND2_X2 U103 ( .A1(n103), .A2(n96), .ZN(n94) );
  NAND2_X2 U107 ( .A1(n96), .A2(n99), .ZN(n11) );
  NAND2_X2 U110 ( .A1(A[10]), .A2(B[10]), .ZN(n99) );
  XNOR2_X2 U111 ( .A(n111), .B(n12), .ZN(SUM[9]) );
  NAND2_X2 U121 ( .A1(n168), .A2(n110), .ZN(n12) );
  NAND2_X2 U124 ( .A1(A[9]), .A2(B[9]), .ZN(n110) );
  XOR2_X2 U125 ( .A(n13), .B(n114), .Z(SUM[8]) );
  NAND2_X2 U127 ( .A1(n169), .A2(n113), .ZN(n13) );
  NAND2_X2 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n113) );
  XOR2_X2 U131 ( .A(n14), .B(n122), .Z(SUM[7]) );
  NAND2_X2 U134 ( .A1(n130), .A2(n118), .ZN(n116) );
  NAND2_X2 U138 ( .A1(n170), .A2(n121), .ZN(n14) );
  NAND2_X2 U141 ( .A1(A[7]), .A2(B[7]), .ZN(n121) );
  XOR2_X2 U142 ( .A(n15), .B(n129), .Z(SUM[6]) );
  NAND2_X2 U148 ( .A1(n171), .A2(n128), .ZN(n15) );
  NAND2_X2 U151 ( .A1(A[6]), .A2(B[6]), .ZN(n128) );
  XOR2_X2 U152 ( .A(n16), .B(n138), .Z(SUM[5]) );
  NAND2_X2 U160 ( .A1(n172), .A2(n137), .ZN(n16) );
  NAND2_X2 U163 ( .A1(A[5]), .A2(B[5]), .ZN(n137) );
  XNOR2_X2 U164 ( .A(n143), .B(n17), .ZN(SUM[4]) );
  NAND2_X2 U168 ( .A1(n173), .A2(n142), .ZN(n17) );
  NAND2_X2 U171 ( .A1(A[4]), .A2(B[4]), .ZN(n142) );
  XNOR2_X2 U172 ( .A(n149), .B(n18), .ZN(SUM[3]) );
  NAND2_X2 U177 ( .A1(n174), .A2(n148), .ZN(n18) );
  NAND2_X2 U180 ( .A1(A[3]), .A2(B[3]), .ZN(n148) );
  XOR2_X2 U181 ( .A(n19), .B(n152), .Z(SUM[2]) );
  NAND2_X2 U183 ( .A1(n175), .A2(n151), .ZN(n19) );
  NAND2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n151) );
  XOR2_X2 U187 ( .A(n157), .B(n20), .Z(SUM[1]) );
  NAND2_X2 U190 ( .A1(n176), .A2(n155), .ZN(n20) );
  NAND2_X2 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n155) );
  NAND2_X2 U198 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  OR2_X4 U202 ( .A1(n30), .A2(n27), .ZN(n247) );
  AND2_X1 U203 ( .A1(n249), .A2(n157), .ZN(SUM[0]) );
  NOR2_X1 U204 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  NOR2_X1 U205 ( .A1(A[18]), .A2(B[18]), .ZN(n34) );
  OAI21_X1 U206 ( .B1(n114), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X1 U207 ( .B1(n86), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U208 ( .B1(n114), .B2(n56), .A(n57), .ZN(n55) );
  AOI21_X4 U209 ( .B1(n115), .B2(n47), .A(n48), .ZN(n1) );
  AOI21_X1 U210 ( .B1(n86), .B2(n67), .A(n68), .ZN(n66) );
  AOI21_X1 U211 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U212 ( .B1(n1), .B2(n37), .A(n38), .ZN(n36) );
  INV_X1 U213 ( .A(n40), .ZN(n38) );
  OAI21_X1 U214 ( .B1(n114), .B2(n101), .A(n102), .ZN(n100) );
  INV_X1 U215 ( .A(n104), .ZN(n102) );
  NOR2_X1 U216 ( .A1(n69), .A2(n60), .ZN(n58) );
  OAI21_X1 U217 ( .B1(n133), .B2(n125), .A(n128), .ZN(n124) );
  NOR2_X1 U218 ( .A1(n132), .A2(n125), .ZN(n123) );
  NOR2_X1 U219 ( .A1(n80), .A2(n73), .ZN(n67) );
  OAI21_X1 U220 ( .B1(n114), .B2(n94), .A(n95), .ZN(n93) );
  OAI21_X1 U221 ( .B1(n1), .B2(n44), .A(n45), .ZN(n43) );
  NOR2_X1 U222 ( .A1(n141), .A2(n136), .ZN(n130) );
  NOR2_X1 U223 ( .A1(n112), .A2(n109), .ZN(n103) );
  NOR2_X1 U224 ( .A1(n150), .A2(n147), .ZN(n145) );
  OAI21_X1 U225 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  OAI21_X1 U226 ( .B1(n120), .B2(n128), .A(n121), .ZN(n119) );
  NOR2_X1 U227 ( .A1(n44), .A2(n41), .ZN(n39) );
  NOR2_X1 U228 ( .A1(n98), .A2(n91), .ZN(n89) );
  NOR2_X1 U229 ( .A1(n60), .A2(n53), .ZN(n51) );
  OAI21_X1 U230 ( .B1(n31), .B2(n27), .A(n28), .ZN(n26) );
  NOR2_X1 U231 ( .A1(A[16]), .A2(B[16]), .ZN(n44) );
  NOR2_X1 U232 ( .A1(A[12]), .A2(B[12]), .ZN(n80) );
  NOR2_X1 U233 ( .A1(n83), .A2(n49), .ZN(n47) );
  OAI21_X2 U234 ( .B1(n84), .B2(n49), .A(n50), .ZN(n48) );
  OAI21_X1 U235 ( .B1(n1), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X1 U236 ( .B1(n114), .B2(n83), .A(n84), .ZN(n82) );
  OAI21_X1 U237 ( .B1(n114), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U238 ( .B1(n40), .B2(n32), .A(n33), .ZN(n31) );
  OAI21_X2 U239 ( .B1(n109), .B2(n113), .A(n110), .ZN(n104) );
  AOI21_X2 U240 ( .B1(n145), .B2(n153), .A(n146), .ZN(n144) );
  OAI21_X2 U241 ( .B1(n73), .B2(n81), .A(n74), .ZN(n68) );
  OAI21_X2 U242 ( .B1(n136), .B2(n142), .A(n137), .ZN(n131) );
  OAI21_X2 U243 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI21_X2 U244 ( .B1(n144), .B2(n116), .A(n117), .ZN(n115) );
  AOI21_X2 U245 ( .B1(n118), .B2(n131), .A(n119), .ZN(n117) );
  NOR2_X2 U246 ( .A1(n125), .A2(n120), .ZN(n118) );
  AOI21_X2 U247 ( .B1(n51), .B2(n68), .A(n52), .ZN(n50) );
  OAI21_X2 U248 ( .B1(n53), .B2(n63), .A(n54), .ZN(n52) );
  AOI21_X2 U249 ( .B1(n143), .B2(n123), .A(n124), .ZN(n122) );
  AOI21_X2 U250 ( .B1(n143), .B2(n173), .A(n140), .ZN(n138) );
  OAI21_X2 U251 ( .B1(n154), .B2(n157), .A(n155), .ZN(n153) );
  AOI21_X2 U252 ( .B1(n89), .B2(n104), .A(n90), .ZN(n84) );
  OAI21_X2 U253 ( .B1(n91), .B2(n99), .A(n92), .ZN(n90) );
  OAI21_X1 U254 ( .B1(n70), .B2(n60), .A(n63), .ZN(n59) );
  AOI21_X2 U255 ( .B1(n86), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X1 U256 ( .B1(n104), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U257 ( .B1(n114), .B2(n112), .A(n113), .ZN(n111) );
  OAI21_X1 U258 ( .B1(n152), .B2(n150), .A(n151), .ZN(n149) );
  NOR2_X2 U259 ( .A1(A[14]), .A2(B[14]), .ZN(n60) );
  NOR2_X2 U260 ( .A1(A[6]), .A2(B[6]), .ZN(n125) );
  NOR2_X2 U261 ( .A1(A[13]), .A2(B[13]), .ZN(n73) );
  NOR2_X2 U262 ( .A1(A[15]), .A2(B[15]), .ZN(n53) );
  NOR2_X2 U263 ( .A1(A[11]), .A2(B[11]), .ZN(n91) );
  NOR2_X2 U264 ( .A1(A[9]), .A2(B[9]), .ZN(n109) );
  NOR2_X2 U265 ( .A1(A[5]), .A2(B[5]), .ZN(n136) );
  NOR2_X2 U266 ( .A1(A[7]), .A2(B[7]), .ZN(n120) );
  NOR2_X2 U267 ( .A1(A[17]), .A2(B[17]), .ZN(n41) );
  NOR2_X2 U268 ( .A1(A[3]), .A2(B[3]), .ZN(n147) );
  NOR2_X2 U269 ( .A1(A[19]), .A2(B[19]), .ZN(n27) );
  NOR2_X1 U270 ( .A1(A[8]), .A2(B[8]), .ZN(n112) );
  NOR2_X2 U271 ( .A1(A[1]), .A2(B[1]), .ZN(n154) );
  NOR2_X1 U272 ( .A1(A[10]), .A2(B[10]), .ZN(n98) );
  NOR2_X1 U273 ( .A1(A[4]), .A2(B[4]), .ZN(n141) );
  OAI21_X2 U274 ( .B1(n1), .B2(n247), .A(n24), .ZN(SUM[20]) );
  OR2_X1 U275 ( .A1(A[0]), .A2(B[0]), .ZN(n249) );
  INV_X4 U276 ( .A(n99), .ZN(n97) );
  INV_X4 U277 ( .A(n84), .ZN(n86) );
  INV_X4 U278 ( .A(n83), .ZN(n85) );
  INV_X4 U279 ( .A(n81), .ZN(n79) );
  INV_X4 U280 ( .A(n68), .ZN(n70) );
  INV_X4 U281 ( .A(n67), .ZN(n69) );
  INV_X4 U282 ( .A(n39), .ZN(n37) );
  INV_X4 U283 ( .A(n35), .ZN(n33) );
  INV_X4 U284 ( .A(n26), .ZN(n24) );
  INV_X4 U285 ( .A(n154), .ZN(n176) );
  INV_X4 U286 ( .A(n150), .ZN(n175) );
  INV_X4 U287 ( .A(n147), .ZN(n174) );
  INV_X4 U288 ( .A(n136), .ZN(n172) );
  INV_X4 U289 ( .A(n125), .ZN(n171) );
  INV_X4 U290 ( .A(n120), .ZN(n170) );
  INV_X4 U291 ( .A(n112), .ZN(n169) );
  INV_X4 U292 ( .A(n109), .ZN(n168) );
  INV_X4 U293 ( .A(n98), .ZN(n96) );
  INV_X4 U294 ( .A(n91), .ZN(n166) );
  INV_X4 U295 ( .A(n80), .ZN(n78) );
  INV_X4 U296 ( .A(n73), .ZN(n164) );
  INV_X4 U297 ( .A(n60), .ZN(n163) );
  INV_X4 U298 ( .A(n53), .ZN(n162) );
  INV_X4 U299 ( .A(n44), .ZN(n161) );
  INV_X4 U300 ( .A(n41), .ZN(n160) );
  INV_X4 U301 ( .A(n34), .ZN(n32) );
  INV_X4 U302 ( .A(n27), .ZN(n158) );
  INV_X4 U303 ( .A(n153), .ZN(n152) );
  INV_X4 U304 ( .A(n144), .ZN(n143) );
  INV_X4 U305 ( .A(n142), .ZN(n140) );
  INV_X4 U306 ( .A(n141), .ZN(n173) );
  INV_X4 U307 ( .A(n131), .ZN(n133) );
  INV_X4 U308 ( .A(n130), .ZN(n132) );
  INV_X4 U309 ( .A(n115), .ZN(n114) );
  INV_X4 U310 ( .A(n103), .ZN(n101) );
endmodule


module pipleline_stage_3 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n106;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;

  pipleline_stage_3_DW01_add_1 add_268 ( .A({1'b0, divided[26:7]}), .B({1'b0, 
        divisor}), .CI(1'b0), .SUM(stage_result) );
  BUF_X4 U5 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U6 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U7 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U8 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U9 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U10 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U11 ( .A(divided[0]), .Z(stage_out[1]) );
  INV_X16 U12 ( .A(n106), .ZN(q) );
  XNOR2_X2 U13 ( .A(divided[27]), .B(stage_result[20]), .ZN(n106) );
  MUX2_X2 U14 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U15 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U16 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U17 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U18 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U19 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U20 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U21 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U22 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U23 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U24 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U25 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U26 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U27 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U28 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U29 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U30 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U31 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U32 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U33 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n24, n26, n27, n28, n29, n30, n31, n33, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64, n65, n66, n67,
         n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n128, n129, n130, n131, n132, n133, n136, n137, n138, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n157, n158, n160, n161, n162, n163, n164, n166,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n247, n248,
         n250;

  XNOR2_X2 U3 ( .A(n29), .B(n2), .ZN(SUM[19]) );
  NAND2_X2 U9 ( .A1(n158), .A2(n28), .ZN(n2) );
  NAND2_X2 U12 ( .A1(A[19]), .A2(B[19]), .ZN(n28) );
  XNOR2_X2 U13 ( .A(n36), .B(n3), .ZN(SUM[18]) );
  NAND2_X2 U15 ( .A1(n39), .A2(n247), .ZN(n30) );
  NAND2_X2 U19 ( .A1(n247), .A2(n35), .ZN(n3) );
  NAND2_X2 U22 ( .A1(A[18]), .A2(B[18]), .ZN(n35) );
  XNOR2_X2 U23 ( .A(n43), .B(n4), .ZN(SUM[17]) );
  NAND2_X2 U29 ( .A1(n160), .A2(n42), .ZN(n4) );
  NAND2_X2 U32 ( .A1(A[17]), .A2(B[17]), .ZN(n42) );
  XOR2_X2 U33 ( .A(n5), .B(n1), .Z(SUM[16]) );
  NAND2_X2 U35 ( .A1(n161), .A2(n45), .ZN(n5) );
  NAND2_X2 U38 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U39 ( .A(n55), .B(n6), .ZN(SUM[15]) );
  NAND2_X2 U43 ( .A1(n67), .A2(n51), .ZN(n49) );
  NAND2_X2 U47 ( .A1(n162), .A2(n54), .ZN(n6) );
  NAND2_X2 U50 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  XNOR2_X2 U51 ( .A(n64), .B(n7), .ZN(SUM[14]) );
  NAND2_X2 U53 ( .A1(n58), .A2(n85), .ZN(n56) );
  NAND2_X2 U59 ( .A1(n163), .A2(n63), .ZN(n7) );
  NAND2_X2 U62 ( .A1(A[14]), .A2(B[14]), .ZN(n63) );
  XNOR2_X2 U63 ( .A(n75), .B(n8), .ZN(SUM[13]) );
  NAND2_X2 U65 ( .A1(n85), .A2(n67), .ZN(n65) );
  NAND2_X2 U73 ( .A1(n164), .A2(n74), .ZN(n8) );
  NAND2_X2 U76 ( .A1(A[13]), .A2(B[13]), .ZN(n74) );
  XNOR2_X2 U77 ( .A(n82), .B(n9), .ZN(SUM[12]) );
  NAND2_X2 U79 ( .A1(n85), .A2(n78), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n78), .A2(n81), .ZN(n9) );
  NAND2_X2 U86 ( .A1(A[12]), .A2(B[12]), .ZN(n81) );
  XNOR2_X2 U87 ( .A(n93), .B(n10), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(n103), .A2(n89), .ZN(n83) );
  NAND2_X2 U97 ( .A1(n166), .A2(n92), .ZN(n10) );
  NAND2_X2 U100 ( .A1(A[11]), .A2(B[11]), .ZN(n92) );
  XNOR2_X2 U101 ( .A(n100), .B(n11), .ZN(SUM[10]) );
  NAND2_X2 U103 ( .A1(n103), .A2(n96), .ZN(n94) );
  NAND2_X2 U107 ( .A1(n96), .A2(n99), .ZN(n11) );
  NAND2_X2 U110 ( .A1(A[10]), .A2(B[10]), .ZN(n99) );
  XNOR2_X2 U111 ( .A(n111), .B(n12), .ZN(SUM[9]) );
  NAND2_X2 U121 ( .A1(n168), .A2(n110), .ZN(n12) );
  NAND2_X2 U124 ( .A1(A[9]), .A2(B[9]), .ZN(n110) );
  XOR2_X2 U125 ( .A(n13), .B(n114), .Z(SUM[8]) );
  NAND2_X2 U127 ( .A1(n169), .A2(n113), .ZN(n13) );
  NAND2_X2 U130 ( .A1(A[8]), .A2(B[8]), .ZN(n113) );
  XOR2_X2 U131 ( .A(n14), .B(n122), .Z(SUM[7]) );
  NAND2_X2 U134 ( .A1(n130), .A2(n118), .ZN(n116) );
  NAND2_X2 U138 ( .A1(n170), .A2(n121), .ZN(n14) );
  NAND2_X2 U141 ( .A1(A[7]), .A2(B[7]), .ZN(n121) );
  XOR2_X2 U142 ( .A(n15), .B(n129), .Z(SUM[6]) );
  NAND2_X2 U148 ( .A1(n171), .A2(n128), .ZN(n15) );
  NAND2_X2 U151 ( .A1(A[6]), .A2(B[6]), .ZN(n128) );
  XOR2_X2 U152 ( .A(n16), .B(n138), .Z(SUM[5]) );
  NAND2_X2 U160 ( .A1(n172), .A2(n137), .ZN(n16) );
  NAND2_X2 U163 ( .A1(A[5]), .A2(B[5]), .ZN(n137) );
  XNOR2_X2 U164 ( .A(n143), .B(n17), .ZN(SUM[4]) );
  NAND2_X2 U168 ( .A1(n173), .A2(n142), .ZN(n17) );
  NAND2_X2 U171 ( .A1(A[4]), .A2(B[4]), .ZN(n142) );
  XNOR2_X2 U172 ( .A(n149), .B(n18), .ZN(SUM[3]) );
  NAND2_X2 U177 ( .A1(n174), .A2(n148), .ZN(n18) );
  NAND2_X2 U180 ( .A1(A[3]), .A2(B[3]), .ZN(n148) );
  XOR2_X2 U181 ( .A(n19), .B(n152), .Z(SUM[2]) );
  NAND2_X2 U183 ( .A1(n175), .A2(n151), .ZN(n19) );
  NAND2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n151) );
  XOR2_X2 U187 ( .A(n157), .B(n20), .Z(SUM[1]) );
  NAND2_X2 U190 ( .A1(n176), .A2(n155), .ZN(n20) );
  NAND2_X2 U193 ( .A1(A[1]), .A2(B[1]), .ZN(n155) );
  NAND2_X2 U198 ( .A1(A[0]), .A2(B[0]), .ZN(n157) );
  OR2_X2 U202 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  OR2_X4 U203 ( .A1(n30), .A2(n27), .ZN(n248) );
  AND2_X1 U204 ( .A1(n250), .A2(n157), .ZN(SUM[0]) );
  NOR2_X1 U205 ( .A1(A[2]), .A2(B[2]), .ZN(n150) );
  OAI21_X1 U206 ( .B1(n114), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X1 U207 ( .B1(n86), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U208 ( .B1(n114), .B2(n56), .A(n57), .ZN(n55) );
  AOI21_X4 U209 ( .B1(n115), .B2(n47), .A(n48), .ZN(n1) );
  AOI21_X1 U210 ( .B1(n86), .B2(n67), .A(n68), .ZN(n66) );
  AOI21_X1 U211 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U212 ( .B1(n1), .B2(n37), .A(n38), .ZN(n36) );
  INV_X1 U213 ( .A(n40), .ZN(n38) );
  OAI21_X1 U214 ( .B1(n114), .B2(n101), .A(n102), .ZN(n100) );
  INV_X1 U215 ( .A(n104), .ZN(n102) );
  NOR2_X1 U216 ( .A1(n69), .A2(n60), .ZN(n58) );
  OAI21_X1 U217 ( .B1(n133), .B2(n125), .A(n128), .ZN(n124) );
  NOR2_X1 U218 ( .A1(n132), .A2(n125), .ZN(n123) );
  NOR2_X1 U219 ( .A1(n80), .A2(n73), .ZN(n67) );
  OAI21_X1 U220 ( .B1(n114), .B2(n94), .A(n95), .ZN(n93) );
  OAI21_X1 U221 ( .B1(n1), .B2(n44), .A(n45), .ZN(n43) );
  NOR2_X1 U222 ( .A1(n141), .A2(n136), .ZN(n130) );
  NOR2_X1 U223 ( .A1(n112), .A2(n109), .ZN(n103) );
  NOR2_X1 U224 ( .A1(n150), .A2(n147), .ZN(n145) );
  OAI21_X1 U225 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  OAI21_X1 U226 ( .B1(n120), .B2(n128), .A(n121), .ZN(n119) );
  NOR2_X1 U227 ( .A1(n44), .A2(n41), .ZN(n39) );
  NOR2_X1 U228 ( .A1(n98), .A2(n91), .ZN(n89) );
  NOR2_X1 U229 ( .A1(n60), .A2(n53), .ZN(n51) );
  OAI21_X1 U230 ( .B1(n31), .B2(n27), .A(n28), .ZN(n26) );
  NOR2_X1 U231 ( .A1(A[16]), .A2(B[16]), .ZN(n44) );
  NOR2_X1 U232 ( .A1(A[12]), .A2(B[12]), .ZN(n80) );
  NOR2_X1 U233 ( .A1(n83), .A2(n49), .ZN(n47) );
  OAI21_X2 U234 ( .B1(n84), .B2(n49), .A(n50), .ZN(n48) );
  OAI21_X1 U235 ( .B1(n1), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X1 U236 ( .B1(n114), .B2(n83), .A(n84), .ZN(n82) );
  OAI21_X1 U237 ( .B1(n114), .B2(n65), .A(n66), .ZN(n64) );
  AOI21_X1 U238 ( .B1(n40), .B2(n247), .A(n33), .ZN(n31) );
  OAI21_X2 U239 ( .B1(n109), .B2(n113), .A(n110), .ZN(n104) );
  AOI21_X2 U240 ( .B1(n145), .B2(n153), .A(n146), .ZN(n144) );
  OAI21_X2 U241 ( .B1(n73), .B2(n81), .A(n74), .ZN(n68) );
  OAI21_X2 U242 ( .B1(n136), .B2(n142), .A(n137), .ZN(n131) );
  OAI21_X2 U243 ( .B1(n41), .B2(n45), .A(n42), .ZN(n40) );
  OAI21_X2 U244 ( .B1(n144), .B2(n116), .A(n117), .ZN(n115) );
  AOI21_X2 U245 ( .B1(n118), .B2(n131), .A(n119), .ZN(n117) );
  NOR2_X2 U246 ( .A1(n125), .A2(n120), .ZN(n118) );
  AOI21_X2 U247 ( .B1(n51), .B2(n68), .A(n52), .ZN(n50) );
  OAI21_X2 U248 ( .B1(n53), .B2(n63), .A(n54), .ZN(n52) );
  AOI21_X2 U249 ( .B1(n143), .B2(n123), .A(n124), .ZN(n122) );
  AOI21_X2 U250 ( .B1(n143), .B2(n173), .A(n140), .ZN(n138) );
  OAI21_X2 U251 ( .B1(n154), .B2(n157), .A(n155), .ZN(n153) );
  AOI21_X2 U252 ( .B1(n89), .B2(n104), .A(n90), .ZN(n84) );
  OAI21_X2 U253 ( .B1(n91), .B2(n99), .A(n92), .ZN(n90) );
  OAI21_X1 U254 ( .B1(n70), .B2(n60), .A(n63), .ZN(n59) );
  AOI21_X2 U255 ( .B1(n86), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X1 U256 ( .B1(n104), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U257 ( .B1(n114), .B2(n112), .A(n113), .ZN(n111) );
  OAI21_X1 U258 ( .B1(n152), .B2(n150), .A(n151), .ZN(n149) );
  NOR2_X2 U259 ( .A1(A[14]), .A2(B[14]), .ZN(n60) );
  NOR2_X2 U260 ( .A1(A[6]), .A2(B[6]), .ZN(n125) );
  NOR2_X2 U261 ( .A1(A[13]), .A2(B[13]), .ZN(n73) );
  NOR2_X2 U262 ( .A1(A[15]), .A2(B[15]), .ZN(n53) );
  NOR2_X2 U263 ( .A1(A[11]), .A2(B[11]), .ZN(n91) );
  NOR2_X2 U264 ( .A1(A[9]), .A2(B[9]), .ZN(n109) );
  NOR2_X2 U265 ( .A1(A[5]), .A2(B[5]), .ZN(n136) );
  NOR2_X2 U266 ( .A1(A[7]), .A2(B[7]), .ZN(n120) );
  NOR2_X2 U267 ( .A1(A[17]), .A2(B[17]), .ZN(n41) );
  NOR2_X2 U268 ( .A1(A[3]), .A2(B[3]), .ZN(n147) );
  NOR2_X2 U269 ( .A1(A[19]), .A2(B[19]), .ZN(n27) );
  NOR2_X1 U270 ( .A1(A[8]), .A2(B[8]), .ZN(n112) );
  NOR2_X2 U271 ( .A1(A[1]), .A2(B[1]), .ZN(n154) );
  NOR2_X1 U272 ( .A1(A[10]), .A2(B[10]), .ZN(n98) );
  NOR2_X1 U273 ( .A1(A[4]), .A2(B[4]), .ZN(n141) );
  OAI21_X2 U274 ( .B1(n1), .B2(n248), .A(n24), .ZN(SUM[20]) );
  OR2_X1 U275 ( .A1(A[0]), .A2(B[0]), .ZN(n250) );
  INV_X4 U276 ( .A(n99), .ZN(n97) );
  INV_X4 U277 ( .A(n84), .ZN(n86) );
  INV_X4 U278 ( .A(n83), .ZN(n85) );
  INV_X4 U279 ( .A(n81), .ZN(n79) );
  INV_X4 U280 ( .A(n68), .ZN(n70) );
  INV_X4 U281 ( .A(n67), .ZN(n69) );
  INV_X4 U282 ( .A(n39), .ZN(n37) );
  INV_X4 U283 ( .A(n35), .ZN(n33) );
  INV_X4 U284 ( .A(n26), .ZN(n24) );
  INV_X4 U285 ( .A(n154), .ZN(n176) );
  INV_X4 U286 ( .A(n150), .ZN(n175) );
  INV_X4 U287 ( .A(n147), .ZN(n174) );
  INV_X4 U288 ( .A(n136), .ZN(n172) );
  INV_X4 U289 ( .A(n125), .ZN(n171) );
  INV_X4 U290 ( .A(n120), .ZN(n170) );
  INV_X4 U291 ( .A(n112), .ZN(n169) );
  INV_X4 U292 ( .A(n109), .ZN(n168) );
  INV_X4 U293 ( .A(n98), .ZN(n96) );
  INV_X4 U294 ( .A(n91), .ZN(n166) );
  INV_X4 U295 ( .A(n80), .ZN(n78) );
  INV_X4 U296 ( .A(n73), .ZN(n164) );
  INV_X4 U297 ( .A(n60), .ZN(n163) );
  INV_X4 U298 ( .A(n53), .ZN(n162) );
  INV_X4 U299 ( .A(n44), .ZN(n161) );
  INV_X4 U300 ( .A(n41), .ZN(n160) );
  INV_X4 U301 ( .A(n27), .ZN(n158) );
  INV_X4 U302 ( .A(n153), .ZN(n152) );
  INV_X4 U303 ( .A(n144), .ZN(n143) );
  INV_X4 U304 ( .A(n142), .ZN(n140) );
  INV_X4 U305 ( .A(n141), .ZN(n173) );
  INV_X4 U306 ( .A(n131), .ZN(n133) );
  INV_X4 U307 ( .A(n130), .ZN(n132) );
  INV_X4 U308 ( .A(n115), .ZN(n114) );
  INV_X4 U309 ( .A(n103), .ZN(n101) );
endmodule


module pipleline_stage_2 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n106;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;

  pipleline_stage_2_DW01_add_1 add_268 ( .A({1'b0, divided[26:7]}), .B({1'b0, 
        divisor}), .CI(1'b0), .SUM(stage_result) );
  BUF_X4 U5 ( .A(divided[0]), .Z(stage_out[1]) );
  BUF_X4 U6 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U7 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U8 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U9 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U10 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U11 ( .A(divided[6]), .Z(stage_out[7]) );
  INV_X16 U12 ( .A(n106), .ZN(q) );
  XNOR2_X2 U13 ( .A(divided[27]), .B(stage_result[20]), .ZN(n106) );
  MUX2_X2 U14 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U15 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U16 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U17 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U18 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U19 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U20 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U21 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U22 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U23 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U24 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U25 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U26 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U27 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U28 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U29 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U30 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U31 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U32 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U33 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_0 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   U3_DATA1_0, U3_DATA1_1, U3_DATA1_2, U3_DATA1_3, U3_DATA1_4,
         U3_DATA1_5, U3_DATA1_6, U3_DATA1_7, U3_DATA1_8, U3_DATA1_9,
         U3_DATA1_10, U3_DATA1_11, U3_DATA1_12, U3_DATA1_13, U3_DATA1_14,
         U3_DATA1_15, U3_DATA1_16, U3_DATA1_17, U3_DATA1_18, U3_DATA1_19, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n99, n100, n109;
  wire   [20:2] add_268_carry;
  assign stage_out[0] = 1'b0;

  FA_X1 add_268_U1_1 ( .A(divided[8]), .B(divisor[1]), .CI(n99), .CO(
        add_268_carry[2]), .S(U3_DATA1_1) );
  FA_X1 add_268_U1_2 ( .A(divided[9]), .B(divisor[2]), .CI(add_268_carry[2]), 
        .CO(add_268_carry[3]), .S(U3_DATA1_2) );
  FA_X1 add_268_U1_3 ( .A(divided[10]), .B(divisor[3]), .CI(add_268_carry[3]), 
        .CO(add_268_carry[4]), .S(U3_DATA1_3) );
  FA_X1 add_268_U1_4 ( .A(divided[11]), .B(divisor[4]), .CI(add_268_carry[4]), 
        .CO(add_268_carry[5]), .S(U3_DATA1_4) );
  FA_X1 add_268_U1_5 ( .A(divided[12]), .B(divisor[5]), .CI(add_268_carry[5]), 
        .CO(add_268_carry[6]), .S(U3_DATA1_5) );
  FA_X1 add_268_U1_6 ( .A(divided[13]), .B(divisor[6]), .CI(add_268_carry[6]), 
        .CO(add_268_carry[7]), .S(U3_DATA1_6) );
  FA_X1 add_268_U1_7 ( .A(divided[14]), .B(divisor[7]), .CI(add_268_carry[7]), 
        .CO(add_268_carry[8]), .S(U3_DATA1_7) );
  FA_X1 add_268_U1_8 ( .A(divided[15]), .B(divisor[8]), .CI(add_268_carry[8]), 
        .CO(add_268_carry[9]), .S(U3_DATA1_8) );
  FA_X1 add_268_U1_9 ( .A(divided[16]), .B(divisor[9]), .CI(add_268_carry[9]), 
        .CO(add_268_carry[10]), .S(U3_DATA1_9) );
  FA_X1 add_268_U1_10 ( .A(divided[17]), .B(divisor[10]), .CI(
        add_268_carry[10]), .CO(add_268_carry[11]), .S(U3_DATA1_10) );
  FA_X1 add_268_U1_11 ( .A(divided[18]), .B(divisor[11]), .CI(
        add_268_carry[11]), .CO(add_268_carry[12]), .S(U3_DATA1_11) );
  FA_X1 add_268_U1_12 ( .A(divided[19]), .B(divisor[12]), .CI(
        add_268_carry[12]), .CO(add_268_carry[13]), .S(U3_DATA1_12) );
  FA_X1 add_268_U1_13 ( .A(divided[20]), .B(divisor[13]), .CI(
        add_268_carry[13]), .CO(add_268_carry[14]), .S(U3_DATA1_13) );
  FA_X1 add_268_U1_14 ( .A(divided[21]), .B(divisor[14]), .CI(
        add_268_carry[14]), .CO(add_268_carry[15]), .S(U3_DATA1_14) );
  FA_X1 add_268_U1_15 ( .A(divided[22]), .B(divisor[15]), .CI(
        add_268_carry[15]), .CO(add_268_carry[16]), .S(U3_DATA1_15) );
  FA_X1 add_268_U1_16 ( .A(divided[23]), .B(divisor[16]), .CI(
        add_268_carry[16]), .CO(add_268_carry[17]), .S(U3_DATA1_16) );
  FA_X1 add_268_U1_17 ( .A(divided[24]), .B(divisor[17]), .CI(
        add_268_carry[17]), .CO(add_268_carry[18]), .S(U3_DATA1_17) );
  FA_X1 add_268_U1_18 ( .A(divided[25]), .B(divisor[18]), .CI(
        add_268_carry[18]), .CO(add_268_carry[19]), .S(U3_DATA1_18) );
  FA_X1 add_268_U1_19 ( .A(divided[26]), .B(divisor[19]), .CI(
        add_268_carry[19]), .CO(add_268_carry[20]), .S(U3_DATA1_19) );
  INV_X4 U2 ( .A(n24), .ZN(stage_out[17]) );
  INV_X4 U5 ( .A(n26), .ZN(stage_out[16]) );
  INV_X4 U7 ( .A(n27), .ZN(stage_out[15]) );
  INV_X4 U9 ( .A(n28), .ZN(stage_out[14]) );
  INV_X4 U11 ( .A(n29), .ZN(stage_out[13]) );
  INV_X4 U13 ( .A(n30), .ZN(stage_out[12]) );
  INV_X4 U15 ( .A(n31), .ZN(stage_out[11]) );
  INV_X4 U17 ( .A(n32), .ZN(stage_out[10]) );
  INV_X4 U19 ( .A(n33), .ZN(stage_out[27]) );
  INV_X4 U21 ( .A(n34), .ZN(stage_out[26]) );
  INV_X4 U23 ( .A(n35), .ZN(stage_out[25]) );
  INV_X4 U25 ( .A(n36), .ZN(stage_out[24]) );
  INV_X4 U27 ( .A(n37), .ZN(stage_out[23]) );
  INV_X4 U29 ( .A(n38), .ZN(stage_out[22]) );
  INV_X4 U31 ( .A(n39), .ZN(stage_out[21]) );
  INV_X4 U33 ( .A(n40), .ZN(stage_out[20]) );
  INV_X4 U35 ( .A(n41), .ZN(stage_out[19]) );
  INV_X4 U37 ( .A(n42), .ZN(stage_out[18]) );
  INV_X4 U39 ( .A(n43), .ZN(stage_out[9]) );
  INV_X4 U41 ( .A(n44), .ZN(stage_out[8]) );
  XNOR2_X2 U44 ( .A(divided[27]), .B(add_268_carry[20]), .ZN(n25) );
  AND2_X4 U6 ( .A1(divisor[0]), .A2(divided[7]), .ZN(n99) );
  BUF_X4 U8 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U10 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U12 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U14 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U16 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U18 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U20 ( .A(divided[0]), .Z(stage_out[1]) );
  AOI22_X2 U22 ( .A1(divided[7]), .A2(n25), .B1(U3_DATA1_0), .B2(n100), .ZN(
        n44) );
  AOI22_X2 U24 ( .A1(divided[8]), .A2(n25), .B1(U3_DATA1_1), .B2(n100), .ZN(
        n43) );
  AOI22_X2 U26 ( .A1(divided[17]), .A2(n25), .B1(U3_DATA1_10), .B2(n100), .ZN(
        n42) );
  AOI22_X2 U28 ( .A1(divided[18]), .A2(n25), .B1(U3_DATA1_11), .B2(q), .ZN(n41) );
  AOI22_X2 U30 ( .A1(divided[19]), .A2(n25), .B1(U3_DATA1_12), .B2(n100), .ZN(
        n40) );
  AOI22_X2 U32 ( .A1(divided[20]), .A2(n25), .B1(U3_DATA1_13), .B2(q), .ZN(n39) );
  AOI22_X2 U34 ( .A1(divided[21]), .A2(n25), .B1(U3_DATA1_14), .B2(n100), .ZN(
        n38) );
  AOI22_X2 U36 ( .A1(divided[22]), .A2(n25), .B1(U3_DATA1_15), .B2(q), .ZN(n37) );
  AOI22_X2 U38 ( .A1(divided[23]), .A2(n25), .B1(U3_DATA1_16), .B2(n100), .ZN(
        n36) );
  AOI22_X2 U40 ( .A1(divided[24]), .A2(n25), .B1(U3_DATA1_17), .B2(q), .ZN(n35) );
  AOI22_X2 U42 ( .A1(divided[25]), .A2(n25), .B1(U3_DATA1_18), .B2(n100), .ZN(
        n34) );
  AOI22_X2 U43 ( .A1(divided[26]), .A2(n25), .B1(U3_DATA1_19), .B2(q), .ZN(n33) );
  AOI22_X2 U45 ( .A1(divided[9]), .A2(n25), .B1(U3_DATA1_2), .B2(n100), .ZN(
        n32) );
  AOI22_X2 U46 ( .A1(divided[10]), .A2(n25), .B1(U3_DATA1_3), .B2(q), .ZN(n31)
         );
  AOI22_X2 U47 ( .A1(divided[11]), .A2(n25), .B1(U3_DATA1_4), .B2(n100), .ZN(
        n30) );
  AOI22_X2 U48 ( .A1(divided[12]), .A2(n25), .B1(U3_DATA1_5), .B2(n100), .ZN(
        n29) );
  AOI22_X2 U49 ( .A1(divided[13]), .A2(n25), .B1(U3_DATA1_6), .B2(q), .ZN(n28)
         );
  AOI22_X2 U50 ( .A1(divided[14]), .A2(n25), .B1(U3_DATA1_7), .B2(n100), .ZN(
        n27) );
  AOI22_X2 U51 ( .A1(divided[15]), .A2(n25), .B1(U3_DATA1_8), .B2(q), .ZN(n26)
         );
  AOI22_X2 U52 ( .A1(divided[16]), .A2(n25), .B1(U3_DATA1_9), .B2(n100), .ZN(
        n24) );
  XOR2_X2 U53 ( .A(divided[27]), .B(add_268_carry[20]), .Z(n100) );
  XOR2_X2 U54 ( .A(divided[27]), .B(add_268_carry[20]), .Z(q) );
  INV_X4 U55 ( .A(divided[7]), .ZN(n109) );
  XNOR2_X2 U56 ( .A(divisor[0]), .B(n109), .ZN(U3_DATA1_0) );
endmodule


module pipeline_divider ( clock, reset_n, start, divided, divisor, q, StartOut
 );
  input [27:0] divided;
  input [19:0] divisor;
  output [7:0] q;
  input clock, reset_n, start;
  output StartOut;
  wire   n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n217, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n355, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n491, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n625, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n887, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, U24_Z_1, U24_Z_2, U24_Z_3,
         U24_Z_4, U24_Z_5, U24_Z_6, U24_Z_7, U24_Z_8, U24_Z_9, U24_Z_10,
         U24_Z_11, U24_Z_12, U24_Z_13, U24_Z_14, U24_Z_15, U24_Z_16, U24_Z_17,
         U24_Z_18, U24_Z_19, U24_Z_20, U24_Z_21, U24_Z_22, U24_Z_23, U24_Z_24,
         U24_Z_25, U24_Z_26, U24_Z_27, U24_DATA1_1, U24_DATA1_2, U24_DATA1_3,
         U24_DATA1_4, U24_DATA1_5, U24_DATA1_6, U24_DATA1_7, U24_DATA1_8,
         U24_DATA1_9, U24_DATA1_10, U24_DATA1_11, U24_DATA1_12, U24_DATA1_13,
         U24_DATA1_14, U24_DATA1_15, U24_DATA1_16, U24_DATA1_17, U24_DATA1_18,
         U24_DATA1_19, U24_DATA1_20, U24_DATA1_21, U24_DATA1_22, U24_DATA1_23,
         U24_DATA1_24, U24_DATA1_25, U24_DATA1_26, U24_DATA1_27, U22_Z_0,
         U22_DATA1_0, U21_Z_1, U21_Z_2, U21_Z_3, U21_Z_4, U21_Z_5, U21_Z_6,
         U21_Z_7, U21_Z_8, U21_Z_9, U21_Z_10, U21_Z_11, U21_Z_12, U21_Z_13,
         U21_Z_14, U21_Z_15, U21_Z_16, U21_Z_17, U21_Z_18, U21_Z_19, U21_Z_20,
         U21_Z_21, U21_Z_22, U21_Z_23, U21_Z_24, U21_Z_25, U21_Z_26, U21_Z_27,
         U21_DATA1_1, U21_DATA1_2, U21_DATA1_3, U21_DATA1_4, U21_DATA1_5,
         U21_DATA1_6, U21_DATA1_7, U21_DATA1_8, U21_DATA1_9, U21_DATA1_10,
         U21_DATA1_11, U21_DATA1_12, U21_DATA1_13, U21_DATA1_14, U21_DATA1_15,
         U21_DATA1_16, U21_DATA1_17, U21_DATA1_18, U21_DATA1_19, U21_DATA1_20,
         U21_DATA1_21, U21_DATA1_22, U21_DATA1_23, U21_DATA1_24, U21_DATA1_25,
         U21_DATA1_26, U21_DATA1_27, U20_Z_0, U20_Z_1, U20_Z_2, U20_Z_3,
         U20_Z_4, U20_Z_5, U20_Z_6, U20_Z_7, U20_Z_8, U20_Z_9, U20_Z_10,
         U20_Z_11, U20_Z_12, U20_Z_13, U20_Z_14, U20_Z_15, U20_Z_16, U20_Z_17,
         U20_Z_18, U20_Z_19, U20_DATA1_0, U20_DATA1_1, U20_DATA1_2,
         U20_DATA1_3, U20_DATA1_4, U20_DATA1_5, U20_DATA1_6, U20_DATA1_7,
         U20_DATA1_8, U20_DATA1_9, U20_DATA1_10, U20_DATA1_11, U20_DATA1_12,
         U20_DATA1_13, U20_DATA1_14, U20_DATA1_15, U20_DATA1_16, U20_DATA1_17,
         U20_DATA1_18, U20_DATA1_19, U19_Z_0, U19_Z_1, U19_DATA1_0,
         U19_DATA1_1, U18_Z_1, U18_Z_2, U18_Z_3, U18_Z_4, U18_Z_5, U18_Z_6,
         U18_Z_7, U18_Z_8, U18_Z_9, U18_Z_10, U18_Z_11, U18_Z_12, U18_Z_13,
         U18_Z_14, U18_Z_15, U18_Z_16, U18_Z_17, U18_Z_18, U18_Z_19, U18_Z_20,
         U18_Z_21, U18_Z_22, U18_Z_23, U18_Z_24, U18_Z_25, U18_Z_26, U18_Z_27,
         U18_DATA1_1, U18_DATA1_2, U18_DATA1_3, U18_DATA1_4, U18_DATA1_5,
         U18_DATA1_6, U18_DATA1_7, U18_DATA1_8, U18_DATA1_9, U18_DATA1_10,
         U18_DATA1_11, U18_DATA1_12, U18_DATA1_13, U18_DATA1_14, U18_DATA1_15,
         U18_DATA1_16, U18_DATA1_17, U18_DATA1_18, U18_DATA1_19, U18_DATA1_20,
         U18_DATA1_21, U18_DATA1_22, U18_DATA1_23, U18_DATA1_24, U18_DATA1_25,
         U18_DATA1_26, U18_DATA1_27, U17_Z_0, U17_Z_1, U17_Z_2, U17_Z_3,
         U17_Z_4, U17_Z_5, U17_Z_6, U17_Z_7, U17_Z_8, U17_Z_9, U17_Z_10,
         U17_Z_11, U17_Z_12, U17_Z_13, U17_Z_14, U17_Z_15, U17_Z_16, U17_Z_17,
         U17_Z_18, U17_Z_19, U17_DATA1_0, U17_DATA1_1, U17_DATA1_2,
         U17_DATA1_3, U17_DATA1_4, U17_DATA1_5, U17_DATA1_6, U17_DATA1_7,
         U17_DATA1_8, U17_DATA1_9, U17_DATA1_10, U17_DATA1_11, U17_DATA1_12,
         U17_DATA1_13, U17_DATA1_14, U17_DATA1_15, U17_DATA1_16, U17_DATA1_17,
         U17_DATA1_18, U17_DATA1_19, U16_Z_0, U16_Z_1, U16_Z_2, U16_DATA1_0,
         U16_DATA1_1, U16_DATA1_2, U15_Z_1, U15_Z_2, U15_Z_3, U15_Z_4, U15_Z_5,
         U15_Z_6, U15_Z_7, U15_Z_8, U15_Z_9, U15_Z_10, U15_Z_11, U15_Z_12,
         U15_Z_13, U15_Z_14, U15_Z_15, U15_Z_16, U15_Z_17, U15_Z_18, U15_Z_19,
         U15_Z_20, U15_Z_21, U15_Z_22, U15_Z_23, U15_Z_24, U15_Z_25, U15_Z_26,
         U15_Z_27, U15_DATA1_1, U15_DATA1_2, U15_DATA1_3, U15_DATA1_4,
         U15_DATA1_5, U15_DATA1_6, U15_DATA1_7, U15_DATA1_8, U15_DATA1_9,
         U15_DATA1_10, U15_DATA1_11, U15_DATA1_12, U15_DATA1_13, U15_DATA1_14,
         U15_DATA1_15, U15_DATA1_16, U15_DATA1_17, U15_DATA1_18, U15_DATA1_19,
         U15_DATA1_20, U15_DATA1_21, U15_DATA1_22, U15_DATA1_23, U15_DATA1_24,
         U15_DATA1_25, U15_DATA1_26, U15_DATA1_27, U14_Z_0, U14_Z_1, U14_Z_2,
         U14_Z_3, U14_Z_4, U14_Z_5, U14_Z_6, U14_Z_7, U14_Z_8, U14_Z_9,
         U14_Z_10, U14_Z_11, U14_Z_12, U14_Z_13, U14_Z_14, U14_Z_15, U14_Z_16,
         U14_Z_17, U14_Z_18, U14_Z_19, U14_DATA1_0, U14_DATA1_1, U14_DATA1_2,
         U14_DATA1_3, U14_DATA1_4, U14_DATA1_5, U14_DATA1_6, U14_DATA1_7,
         U14_DATA1_8, U14_DATA1_9, U14_DATA1_10, U14_DATA1_11, U14_DATA1_12,
         U14_DATA1_13, U14_DATA1_14, U14_DATA1_15, U14_DATA1_16, U14_DATA1_17,
         U14_DATA1_18, U14_DATA1_19, U13_Z_0, U13_Z_1, U13_Z_2, U13_Z_3,
         U13_DATA1_0, U13_DATA1_1, U13_DATA1_2, U13_DATA1_3, U12_Z_1, U12_Z_2,
         U12_Z_3, U12_Z_4, U12_Z_5, U12_Z_6, U12_Z_7, U12_Z_8, U12_Z_9,
         U12_Z_10, U12_Z_11, U12_Z_12, U12_Z_13, U12_Z_14, U12_Z_15, U12_Z_16,
         U12_Z_17, U12_Z_18, U12_Z_19, U12_Z_20, U12_Z_21, U12_Z_22, U12_Z_23,
         U12_Z_24, U12_Z_25, U12_Z_26, U12_Z_27, U12_DATA1_1, U12_DATA1_2,
         U12_DATA1_3, U12_DATA1_4, U12_DATA1_5, U12_DATA1_6, U12_DATA1_7,
         U12_DATA1_8, U12_DATA1_9, U12_DATA1_10, U12_DATA1_11, U12_DATA1_12,
         U12_DATA1_13, U12_DATA1_14, U12_DATA1_15, U12_DATA1_16, U12_DATA1_17,
         U12_DATA1_18, U12_DATA1_19, U12_DATA1_20, U12_DATA1_21, U12_DATA1_22,
         U12_DATA1_23, U12_DATA1_24, U12_DATA1_25, U12_DATA1_26, U12_DATA1_27,
         U11_Z_0, U11_Z_1, U11_Z_2, U11_Z_3, U11_Z_4, U11_Z_5, U11_Z_6,
         U11_Z_7, U11_Z_8, U11_Z_9, U11_Z_10, U11_Z_11, U11_Z_12, U11_Z_13,
         U11_Z_14, U11_Z_15, U11_Z_16, U11_Z_17, U11_Z_18, U11_Z_19,
         U11_DATA1_0, U11_DATA1_1, U11_DATA1_2, U11_DATA1_3, U11_DATA1_4,
         U11_DATA1_5, U11_DATA1_6, U11_DATA1_7, U11_DATA1_8, U11_DATA1_9,
         U11_DATA1_10, U11_DATA1_11, U11_DATA1_12, U11_DATA1_13, U11_DATA1_14,
         U11_DATA1_15, U11_DATA1_16, U11_DATA1_17, U11_DATA1_18, U11_DATA1_19,
         U10_Z_0, U10_Z_1, U10_Z_2, U10_Z_3, U10_Z_4, U10_DATA1_0, U10_DATA1_1,
         U10_DATA1_2, U10_DATA1_3, U10_DATA1_4, U9_Z_1, U9_Z_2, U9_Z_3, U9_Z_4,
         U9_Z_5, U9_Z_6, U9_Z_7, U9_Z_8, U9_Z_9, U9_Z_10, U9_Z_11, U9_Z_12,
         U9_Z_13, U9_Z_14, U9_Z_15, U9_Z_16, U9_Z_17, U9_Z_18, U9_Z_19,
         U9_Z_20, U9_Z_21, U9_Z_22, U9_Z_23, U9_Z_24, U9_Z_25, U9_Z_26,
         U9_Z_27, U9_DATA1_1, U9_DATA1_2, U9_DATA1_3, U9_DATA1_4, U9_DATA1_5,
         U9_DATA1_6, U9_DATA1_7, U9_DATA1_8, U9_DATA1_9, U9_DATA1_10,
         U9_DATA1_11, U9_DATA1_12, U9_DATA1_13, U9_DATA1_14, U9_DATA1_15,
         U9_DATA1_16, U9_DATA1_17, U9_DATA1_18, U9_DATA1_19, U9_DATA1_20,
         U9_DATA1_21, U9_DATA1_22, U9_DATA1_23, U9_DATA1_24, U9_DATA1_25,
         U9_DATA1_26, U9_DATA1_27, U8_Z_0, U8_Z_1, U8_Z_2, U8_Z_3, U8_Z_4,
         U8_Z_5, U8_Z_6, U8_Z_7, U8_Z_8, U8_Z_9, U8_Z_10, U8_Z_11, U8_Z_12,
         U8_Z_13, U8_Z_14, U8_Z_15, U8_Z_16, U8_Z_18, U8_Z_19, U8_DATA1_0,
         U8_DATA1_1, U8_DATA1_2, U8_DATA1_3, U8_DATA1_4, U8_DATA1_5,
         U8_DATA1_6, U8_DATA1_7, U8_DATA1_8, U8_DATA1_9, U8_DATA1_10,
         U8_DATA1_11, U8_DATA1_12, U8_DATA1_13, U8_DATA1_14, U8_DATA1_15,
         U8_DATA1_16, U8_DATA1_17, U8_DATA1_18, U8_DATA1_19, U7_Z_0, U7_Z_1,
         U7_Z_2, U7_Z_3, U7_Z_4, U7_Z_5, U7_DATA1_0, U7_DATA1_1, U7_DATA1_2,
         U7_DATA1_3, U7_DATA1_4, U7_DATA1_5, U6_Z_1, U6_Z_2, U6_Z_3, U6_Z_4,
         U6_Z_5, U6_Z_6, U6_Z_7, U6_Z_8, U6_Z_9, U6_Z_10, U6_Z_11, U6_Z_12,
         U6_Z_13, U6_Z_14, U6_Z_15, U6_Z_16, U6_Z_17, U6_Z_18, U6_Z_19,
         U6_Z_20, U6_Z_21, U6_Z_22, U6_Z_23, U6_Z_24, U6_Z_25, U6_Z_26,
         U6_Z_27, U6_DATA1_1, U6_DATA1_2, U6_DATA1_3, U6_DATA1_4, U6_DATA1_5,
         U6_DATA1_6, U6_DATA1_7, U6_DATA1_8, U6_DATA1_9, U6_DATA1_10,
         U6_DATA1_11, U6_DATA1_12, U6_DATA1_13, U6_DATA1_14, U6_DATA1_15,
         U6_DATA1_16, U6_DATA1_17, U6_DATA1_18, U6_DATA1_19, U6_DATA1_20,
         U6_DATA1_21, U6_DATA1_22, U6_DATA1_23, U6_DATA1_24, U6_DATA1_25,
         U6_DATA1_26, U6_DATA1_27, U5_Z_0, U5_Z_1, U5_Z_2, U5_Z_3, U5_Z_4,
         U5_Z_5, U5_Z_6, U5_Z_7, U5_Z_8, U5_Z_9, U5_Z_10, U5_Z_11, U5_Z_12,
         U5_Z_13, U5_Z_14, U5_Z_15, U5_Z_16, U5_Z_17, U5_Z_18, U5_Z_19,
         U5_DATA1_0, U5_DATA1_1, U5_DATA1_2, U5_DATA1_3, U5_DATA1_4,
         U5_DATA1_5, U5_DATA1_6, U5_DATA1_7, U5_DATA1_8, U5_DATA1_9,
         U5_DATA1_10, U5_DATA1_11, U5_DATA1_12, U5_DATA1_13, U5_DATA1_14,
         U5_DATA1_15, U5_DATA1_16, U5_DATA1_17, U5_DATA1_18, U5_DATA1_19,
         U4_Z_0, U4_Z_1, U4_Z_2, U4_Z_3, U4_Z_4, U4_Z_5, U4_Z_6, U4_DATA1_0,
         U4_DATA1_1, U4_DATA1_2, U4_DATA1_3, U4_DATA1_4, U4_DATA1_5,
         U4_DATA1_6, n21, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1177, n1178, n1179, n1180,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35;
  wire   [104:85] n;

  pipleline_stage_1 stage0 ( .divided(divided), .divisor({n21, n1216, n1217, 
        n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
        n1228, n1229, n1230, n1231, n1232, n1233, n1234}), .q(U22_DATA1_0), 
        .stage_out({U24_DATA1_27, U24_DATA1_26, U24_DATA1_25, U24_DATA1_24, 
        U24_DATA1_23, U24_DATA1_22, U24_DATA1_21, U24_DATA1_20, U24_DATA1_19, 
        U24_DATA1_18, U24_DATA1_17, U24_DATA1_16, U24_DATA1_15, U24_DATA1_14, 
        U24_DATA1_13, U24_DATA1_12, U24_DATA1_11, U24_DATA1_10, U24_DATA1_9, 
        U24_DATA1_8, U24_DATA1_7, U24_DATA1_6, U24_DATA1_5, U24_DATA1_4, 
        U24_DATA1_3, U24_DATA1_2, U24_DATA1_1, SYNOPSYS_UNCONNECTED_1}) );
  pipleline_stage_7 stage1 ( .divided({n936, n935, n934, n933, n932, n931, 
        n930, n929, n928, n927, n926, n925, n924, n923, n922, n921, n920, n919, 
        n918, n917, n916, n915, n914, n913, n912, n911, n910, 1'b0}), 
        .divisor({U20_DATA1_19, U20_DATA1_18, U20_DATA1_17, U20_DATA1_16, 
        U20_DATA1_15, U20_DATA1_14, U20_DATA1_13, U20_DATA1_12, U20_DATA1_11, 
        U20_DATA1_10, U20_DATA1_9, U20_DATA1_8, U20_DATA1_7, U20_DATA1_6, 
        U20_DATA1_5, U20_DATA1_4, U20_DATA1_3, U20_DATA1_2, U20_DATA1_1, 
        U20_DATA1_0}), .q(U19_DATA1_0), .stage_out({U21_DATA1_27, U21_DATA1_26, 
        U21_DATA1_25, U21_DATA1_24, U21_DATA1_23, U21_DATA1_22, U21_DATA1_21, 
        U21_DATA1_20, U21_DATA1_19, U21_DATA1_18, U21_DATA1_17, U21_DATA1_16, 
        U21_DATA1_15, U21_DATA1_14, U21_DATA1_13, U21_DATA1_12, U21_DATA1_11, 
        U21_DATA1_10, U21_DATA1_9, U21_DATA1_8, U21_DATA1_7, U21_DATA1_6, 
        U21_DATA1_5, U21_DATA1_4, U21_DATA1_3, U21_DATA1_2, U21_DATA1_1, 
        SYNOPSYS_UNCONNECTED_2}) );
  pipleline_stage_6 stage2 ( .divided({n807, n806, n805, n804, n803, n802, 
        n801, n800, n799, n798, n797, n796, n795, n794, n793, n792, n791, n790, 
        n789, n788, n787, n786, n785, n784, n783, n782, n781, 1'b0}), 
        .divisor({U17_DATA1_19, U17_DATA1_18, U17_DATA1_17, U17_DATA1_16, 
        U17_DATA1_15, U17_DATA1_14, U17_DATA1_13, U17_DATA1_12, U17_DATA1_11, 
        U17_DATA1_10, U17_DATA1_9, U17_DATA1_8, U17_DATA1_7, U17_DATA1_6, 
        U17_DATA1_5, U17_DATA1_4, U17_DATA1_3, U17_DATA1_2, U17_DATA1_1, 
        U17_DATA1_0}), .q(U16_DATA1_0), .stage_out({U18_DATA1_27, U18_DATA1_26, 
        U18_DATA1_25, U18_DATA1_24, U18_DATA1_23, U18_DATA1_22, U18_DATA1_21, 
        U18_DATA1_20, U18_DATA1_19, U18_DATA1_18, U18_DATA1_17, U18_DATA1_16, 
        U18_DATA1_15, U18_DATA1_14, U18_DATA1_13, U18_DATA1_12, U18_DATA1_11, 
        U18_DATA1_10, U18_DATA1_9, U18_DATA1_8, U18_DATA1_7, U18_DATA1_6, 
        U18_DATA1_5, U18_DATA1_4, U18_DATA1_3, U18_DATA1_2, U18_DATA1_1, 
        SYNOPSYS_UNCONNECTED_3}) );
  pipleline_stage_5 stage3 ( .divided({n676, n675, n674, n673, n672, n671, 
        n670, n669, n668, n667, n666, n665, n664, n663, n662, n661, n660, n659, 
        n658, n657, n656, n655, n654, n653, n652, n651, n650, 1'b0}), 
        .divisor({U14_DATA1_19, U14_DATA1_18, U14_DATA1_17, U14_DATA1_16, 
        U14_DATA1_15, U14_DATA1_14, U14_DATA1_13, U14_DATA1_12, U14_DATA1_11, 
        U14_DATA1_10, U14_DATA1_9, U14_DATA1_8, U14_DATA1_7, U14_DATA1_6, 
        U14_DATA1_5, U14_DATA1_4, U14_DATA1_3, U14_DATA1_2, U14_DATA1_1, 
        U14_DATA1_0}), .q(U13_DATA1_0), .stage_out({U15_DATA1_27, U15_DATA1_26, 
        U15_DATA1_25, U15_DATA1_24, U15_DATA1_23, U15_DATA1_22, U15_DATA1_21, 
        U15_DATA1_20, U15_DATA1_19, U15_DATA1_18, U15_DATA1_17, U15_DATA1_16, 
        U15_DATA1_15, U15_DATA1_14, U15_DATA1_13, U15_DATA1_12, U15_DATA1_11, 
        U15_DATA1_10, U15_DATA1_9, U15_DATA1_8, U15_DATA1_7, U15_DATA1_6, 
        U15_DATA1_5, U15_DATA1_4, U15_DATA1_3, U15_DATA1_2, U15_DATA1_1, 
        SYNOPSYS_UNCONNECTED_4}) );
  pipleline_stage_4 stage4 ( .divided({n543, n542, n541, n540, n539, n538, 
        n537, n536, n535, n534, n533, n532, n531, n530, n529, n528, n527, n526, 
        n525, n524, n523, n522, n521, n520, n519, n518, n517, 1'b0}), 
        .divisor({U11_DATA1_19, U11_DATA1_18, U11_DATA1_17, U11_DATA1_16, 
        U11_DATA1_15, U11_DATA1_14, U11_DATA1_13, U11_DATA1_12, U11_DATA1_11, 
        U11_DATA1_10, U11_DATA1_9, U11_DATA1_8, U11_DATA1_7, U11_DATA1_6, 
        U11_DATA1_5, U11_DATA1_4, U11_DATA1_3, U11_DATA1_2, U11_DATA1_1, 
        U11_DATA1_0}), .q(U10_DATA1_0), .stage_out({U12_DATA1_27, U12_DATA1_26, 
        U12_DATA1_25, U12_DATA1_24, U12_DATA1_23, U12_DATA1_22, U12_DATA1_21, 
        U12_DATA1_20, U12_DATA1_19, U12_DATA1_18, U12_DATA1_17, U12_DATA1_16, 
        U12_DATA1_15, U12_DATA1_14, U12_DATA1_13, U12_DATA1_12, U12_DATA1_11, 
        U12_DATA1_10, U12_DATA1_9, U12_DATA1_8, U12_DATA1_7, U12_DATA1_6, 
        U12_DATA1_5, U12_DATA1_4, U12_DATA1_3, U12_DATA1_2, U12_DATA1_1, 
        SYNOPSYS_UNCONNECTED_5}) );
  pipleline_stage_3 stage5 ( .divided({n408, n407, n406, n405, n404, n403, 
        n402, n401, n400, n399, n398, n397, n396, n395, n394, n393, n392, n391, 
        n390, n389, n388, n387, n386, n385, n384, n383, n382, 1'b0}), 
        .divisor({U8_DATA1_19, U8_DATA1_18, U8_DATA1_17, U8_DATA1_16, 
        U8_DATA1_15, U8_DATA1_14, U8_DATA1_13, U8_DATA1_12, U8_DATA1_11, 
        U8_DATA1_10, U8_DATA1_9, U8_DATA1_8, U8_DATA1_7, U8_DATA1_6, 
        U8_DATA1_5, U8_DATA1_4, U8_DATA1_3, U8_DATA1_2, U8_DATA1_1, U8_DATA1_0}), .q(U7_DATA1_0), .stage_out({U9_DATA1_27, U9_DATA1_26, U9_DATA1_25, 
        U9_DATA1_24, U9_DATA1_23, U9_DATA1_22, U9_DATA1_21, U9_DATA1_20, 
        U9_DATA1_19, U9_DATA1_18, U9_DATA1_17, U9_DATA1_16, U9_DATA1_15, 
        U9_DATA1_14, U9_DATA1_13, U9_DATA1_12, U9_DATA1_11, U9_DATA1_10, 
        U9_DATA1_9, U9_DATA1_8, U9_DATA1_7, U9_DATA1_6, U9_DATA1_5, U9_DATA1_4, 
        U9_DATA1_3, U9_DATA1_2, U9_DATA1_1, SYNOPSYS_UNCONNECTED_6}) );
  pipleline_stage_2 stage6 ( .divided({n271, n270, n269, n268, n267, n266, 
        n265, n264, n263, n262, n261, n260, n259, n258, n257, n256, n255, n254, 
        n253, n252, n251, n250, n249, n248, n247, n246, n245, 1'b0}), 
        .divisor({U5_DATA1_19, U5_DATA1_18, U5_DATA1_17, U5_DATA1_16, 
        U5_DATA1_15, U5_DATA1_14, U5_DATA1_13, U5_DATA1_12, U5_DATA1_11, 
        U5_DATA1_10, U5_DATA1_9, U5_DATA1_8, U5_DATA1_7, U5_DATA1_6, 
        U5_DATA1_5, U5_DATA1_4, U5_DATA1_3, U5_DATA1_2, U5_DATA1_1, U5_DATA1_0}), .q(U4_DATA1_0), .stage_out({U6_DATA1_27, U6_DATA1_26, U6_DATA1_25, 
        U6_DATA1_24, U6_DATA1_23, U6_DATA1_22, U6_DATA1_21, U6_DATA1_20, 
        U6_DATA1_19, U6_DATA1_18, U6_DATA1_17, U6_DATA1_16, U6_DATA1_15, 
        U6_DATA1_14, U6_DATA1_13, U6_DATA1_12, U6_DATA1_11, U6_DATA1_10, 
        U6_DATA1_9, U6_DATA1_8, U6_DATA1_7, U6_DATA1_6, U6_DATA1_5, U6_DATA1_4, 
        U6_DATA1_3, U6_DATA1_2, U6_DATA1_1, SYNOPSYS_UNCONNECTED_7}) );
  pipleline_stage_0 stage7 ( .divided({n132, n131, n130, n129, n128, n127, 
        n126, n125, n124, n123, n122, n121, n120, n119, n118, n117, n116, n115, 
        n114, n113, n112, n111, n110, n109, n108, n107, n106, 1'b0}), 
        .divisor(n), .q(q[0]), .stage_out({SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35}) );
  SDFFR_X2 pipe0_divisor_n_reg_18_ ( .D(1'b0), .SI(start), .SE(n1216), .CK(
        clock), .RN(n1201), .Q(U20_DATA1_18), .QN(n1076) );
  SDFFR_X2 pipe0_divisor_n_reg_17_ ( .D(1'b0), .SI(start), .SE(n1217), .CK(
        clock), .RN(n1203), .Q(U20_DATA1_17), .QN(n1075) );
  SDFFR_X2 pipe0_divisor_n_reg_16_ ( .D(1'b0), .SI(start), .SE(n1218), .CK(
        clock), .RN(n1198), .Q(U20_DATA1_16), .QN(n1083) );
  SDFFR_X2 pipe0_divisor_n_reg_15_ ( .D(1'b0), .SI(start), .SE(n1219), .CK(
        clock), .RN(n1200), .Q(U20_DATA1_15), .QN(n1074) );
  SDFFR_X2 pipe0_divisor_n_reg_14_ ( .D(1'b0), .SI(start), .SE(n1220), .CK(
        clock), .RN(n1201), .Q(U20_DATA1_14), .QN(n1073) );
  SDFFR_X2 pipe0_divisor_n_reg_13_ ( .D(1'b0), .SI(start), .SE(n1221), .CK(
        clock), .RN(n1203), .Q(U20_DATA1_13), .QN(n1072) );
  SDFFR_X2 pipe0_divisor_n_reg_12_ ( .D(1'b0), .SI(start), .SE(n1222), .CK(
        clock), .RN(n1197), .Q(U20_DATA1_12), .QN(n1082) );
  SDFFR_X2 pipe0_divisor_n_reg_10_ ( .D(1'b0), .SI(n1183), .SE(n1224), .CK(
        clock), .RN(n1209), .Q(U20_DATA1_10), .QN(n1081) );
  SDFFR_X2 pipe0_divisor_n_reg_8_ ( .D(1'b0), .SI(n1183), .SE(n1226), .CK(
        clock), .RN(n1191), .Q(U20_DATA1_8), .QN(n1080) );
  SDFFR_X2 pipe0_divisor_n_reg_7_ ( .D(1'b0), .SI(n1183), .SE(n1227), .CK(
        clock), .RN(n1186), .Q(U20_DATA1_7), .QN(n1071) );
  SDFFR_X2 pipe0_divisor_n_reg_6_ ( .D(1'b0), .SI(n1183), .SE(n1228), .CK(
        clock), .RN(n1187), .Q(U20_DATA1_6), .QN(n1070) );
  SDFFR_X2 pipe0_divisor_n_reg_5_ ( .D(1'b0), .SI(n1183), .SE(n1229), .CK(
        clock), .RN(n1192), .Q(U20_DATA1_5), .QN(n1069) );
  SDFFR_X2 pipe0_divisor_n_reg_4_ ( .D(1'b0), .SI(n1183), .SE(n1230), .CK(
        clock), .RN(n1193), .Q(U20_DATA1_4), .QN(n1079) );
  SDFFR_X2 pipe0_divisor_n_reg_2_ ( .D(1'b0), .SI(n1183), .SE(n1232), .CK(
        clock), .RN(n1195), .Q(U20_DATA1_2), .QN(n1078) );
  SDFFR_X2 pipe0_divisor_n_reg_0_ ( .D(1'b0), .SI(n1183), .SE(n1234), .CK(
        clock), .RN(n1196), .Q(U20_DATA1_0), .QN(n1077) );
  DFFR_X1 pipe0_result_reg_26_ ( .D(U24_Z_26), .CK(clock), .RN(n1205), .Q(n935) );
  DFFR_X1 pipe0_result_reg_25_ ( .D(U24_Z_25), .CK(clock), .RN(n1207), .Q(n934) );
  DFFR_X1 pipe0_result_reg_24_ ( .D(U24_Z_24), .CK(clock), .RN(n1208), .Q(n933) );
  DFFR_X1 pipe0_result_reg_23_ ( .D(U24_Z_23), .CK(clock), .RN(n1185), .Q(n932) );
  DFFR_X1 pipe0_result_reg_22_ ( .D(U24_Z_22), .CK(clock), .RN(n1188), .Q(n931) );
  DFFR_X1 pipe0_result_reg_21_ ( .D(U24_Z_21), .CK(clock), .RN(n1190), .Q(n930) );
  DFFR_X1 pipe0_result_reg_20_ ( .D(U24_Z_20), .CK(clock), .RN(n1194), .Q(n929) );
  DFFR_X1 pipe0_result_reg_19_ ( .D(U24_Z_19), .CK(clock), .RN(n1199), .Q(n928) );
  DFFR_X1 pipe0_result_reg_18_ ( .D(U24_Z_18), .CK(clock), .RN(n1202), .Q(n927) );
  DFFR_X1 pipe0_result_reg_17_ ( .D(U24_Z_17), .CK(clock), .RN(n1206), .Q(n926) );
  DFFR_X1 pipe0_result_reg_16_ ( .D(U24_Z_16), .CK(clock), .RN(n1198), .Q(n925) );
  DFFR_X1 pipe0_result_reg_15_ ( .D(U24_Z_15), .CK(clock), .RN(n1200), .Q(n924) );
  DFFR_X1 pipe0_result_reg_14_ ( .D(U24_Z_14), .CK(clock), .RN(n1203), .Q(n923) );
  DFFR_X1 pipe0_result_reg_13_ ( .D(U24_Z_13), .CK(clock), .RN(n1204), .Q(n922) );
  DFFR_X1 pipe0_result_reg_12_ ( .D(U24_Z_12), .CK(clock), .RN(n1205), .Q(n921) );
  DFFR_X1 pipe0_result_reg_11_ ( .D(U24_Z_11), .CK(clock), .RN(n1207), .Q(n920) );
  DFFR_X1 pipe0_result_reg_10_ ( .D(U24_Z_10), .CK(clock), .RN(n1208), .Q(n919) );
  DFFR_X1 pipe0_result_reg_9_ ( .D(U24_Z_9), .CK(clock), .RN(n1185), .Q(n918)
         );
  DFFR_X1 pipe0_result_reg_8_ ( .D(U24_Z_8), .CK(clock), .RN(n1188), .Q(n917)
         );
  DFFR_X1 pipe0_result_reg_7_ ( .D(U24_Z_7), .CK(clock), .RN(n1190), .Q(n916)
         );
  DFFR_X1 pipe1_divisor_n_reg_19_ ( .D(U20_Z_19), .CK(clock), .RN(n1204), .Q(
        U17_DATA1_19) );
  DFFR_X1 pipe1_divisor_n_reg_18_ ( .D(U20_Z_18), .CK(clock), .RN(n1205), .Q(
        U17_DATA1_18), .QN(n1165) );
  DFFR_X1 pipe1_divisor_n_reg_17_ ( .D(U20_Z_17), .CK(clock), .RN(n1207), .Q(
        U17_DATA1_17), .QN(n1124) );
  DFFR_X1 pipe1_divisor_n_reg_15_ ( .D(U20_Z_15), .CK(clock), .RN(n1208), .Q(
        U17_DATA1_15), .QN(n1120) );
  DFFR_X1 pipe1_divisor_n_reg_14_ ( .D(U20_Z_14), .CK(clock), .RN(n1185), .Q(
        U17_DATA1_14), .QN(n1116) );
  DFFR_X1 pipe1_divisor_n_reg_13_ ( .D(U20_Z_13), .CK(clock), .RN(n1188), .Q(
        U17_DATA1_13), .QN(n1112) );
  DFFR_X1 pipe1_divisor_n_reg_12_ ( .D(U20_Z_12), .CK(clock), .RN(n1190), .Q(
        U17_DATA1_12), .QN(n1158) );
  DFFR_X1 pipe1_divisor_n_reg_11_ ( .D(U20_Z_11), .CK(clock), .RN(n1194), .Q(
        U17_DATA1_11), .QN(n1108) );
  DFFR_X1 pipe1_divisor_n_reg_10_ ( .D(U20_Z_10), .CK(clock), .RN(n1202), .Q(
        U17_DATA1_10), .QN(n1154) );
  DFFR_X1 pipe1_divisor_n_reg_9_ ( .D(U20_Z_9), .CK(clock), .RN(n1206), .Q(
        U17_DATA1_9), .QN(n1104) );
  DFFR_X1 pipe1_divisor_n_reg_8_ ( .D(U20_Z_8), .CK(clock), .RN(n1198), .Q(
        U17_DATA1_8), .QN(n1150) );
  DFFR_X1 pipe1_divisor_n_reg_7_ ( .D(U20_Z_7), .CK(clock), .RN(n1200), .Q(
        U17_DATA1_7), .QN(n1100) );
  DFFR_X1 pipe1_divisor_n_reg_6_ ( .D(U20_Z_6), .CK(clock), .RN(n1201), .Q(
        U17_DATA1_6), .QN(n1096) );
  DFFR_X1 pipe1_divisor_n_reg_5_ ( .D(U20_Z_5), .CK(clock), .RN(n1203), .Q(
        U17_DATA1_5), .QN(n1092) );
  DFFR_X1 pipe1_divisor_n_reg_4_ ( .D(U20_Z_4), .CK(clock), .RN(n1204), .Q(
        U17_DATA1_4), .QN(n1146) );
  DFFR_X1 pipe1_divisor_n_reg_3_ ( .D(U20_Z_3), .CK(clock), .RN(n1205), .Q(
        U17_DATA1_3), .QN(n1088) );
  DFFR_X1 pipe1_divisor_n_reg_2_ ( .D(U20_Z_2), .CK(clock), .RN(n1207), .Q(
        U17_DATA1_2), .QN(n1142) );
  DFFR_X1 pipe1_divisor_n_reg_1_ ( .D(U20_Z_1), .CK(clock), .RN(n1208), .Q(
        U17_DATA1_1), .QN(n1084) );
  DFFR_X1 pipe1_divisor_n_reg_0_ ( .D(U20_Z_0), .CK(clock), .RN(n1185), .Q(
        U17_DATA1_0), .QN(n1137) );
  DFFR_X1 pipe1_result_reg_26_ ( .D(U21_Z_26), .CK(clock), .RN(n1190), .Q(n806) );
  DFFR_X1 pipe1_result_reg_25_ ( .D(U21_Z_25), .CK(clock), .RN(n1194), .Q(n805) );
  DFFR_X1 pipe1_result_reg_24_ ( .D(U21_Z_24), .CK(clock), .RN(n1199), .Q(n804) );
  DFFR_X1 pipe1_result_reg_23_ ( .D(U21_Z_23), .CK(clock), .RN(n1202), .Q(n803) );
  DFFR_X1 pipe1_result_reg_22_ ( .D(U21_Z_22), .CK(clock), .RN(n1206), .Q(n802) );
  DFFR_X1 pipe1_result_reg_21_ ( .D(U21_Z_21), .CK(clock), .RN(n1198), .Q(n801) );
  DFFR_X1 pipe1_result_reg_20_ ( .D(U21_Z_20), .CK(clock), .RN(n1200), .Q(n800) );
  DFFR_X1 pipe1_result_reg_19_ ( .D(U21_Z_19), .CK(clock), .RN(n1201), .Q(n799) );
  DFFR_X1 pipe1_result_reg_18_ ( .D(U21_Z_18), .CK(clock), .RN(n1203), .Q(n798) );
  DFFR_X1 pipe1_result_reg_17_ ( .D(U21_Z_17), .CK(clock), .RN(n1205), .Q(n797) );
  DFFR_X1 pipe1_result_reg_16_ ( .D(U21_Z_16), .CK(clock), .RN(n1207), .Q(n796) );
  DFFR_X1 pipe1_result_reg_15_ ( .D(U21_Z_15), .CK(clock), .RN(n1208), .Q(n795) );
  DFFR_X1 pipe1_result_reg_14_ ( .D(U21_Z_14), .CK(clock), .RN(n1185), .Q(n794) );
  DFFR_X1 pipe1_result_reg_13_ ( .D(U21_Z_13), .CK(clock), .RN(n1188), .Q(n793) );
  DFFR_X1 pipe1_result_reg_12_ ( .D(U21_Z_12), .CK(clock), .RN(n1190), .Q(n792) );
  DFFR_X1 pipe1_result_reg_11_ ( .D(U21_Z_11), .CK(clock), .RN(n1194), .Q(n791) );
  DFFR_X1 pipe1_result_reg_10_ ( .D(U21_Z_10), .CK(clock), .RN(n1199), .Q(n790) );
  DFFR_X1 pipe1_result_reg_9_ ( .D(U21_Z_9), .CK(clock), .RN(n1202), .Q(n789)
         );
  DFFR_X1 pipe1_result_reg_8_ ( .D(U21_Z_8), .CK(clock), .RN(n1206), .Q(n788)
         );
  DFFR_X1 pipe1_result_reg_7_ ( .D(U21_Z_7), .CK(clock), .RN(n1198), .Q(n787)
         );
  DFFR_X1 pipe1_result_reg_1_ ( .D(U21_Z_1), .CK(clock), .RN(n1199), .Q(n781)
         );
  DFFR_X1 pipe2_divisor_n_reg_18_ ( .D(U17_Z_18), .CK(clock), .RN(n1202), .Q(
        U14_DATA1_18), .QN(n1166) );
  DFFR_X1 pipe2_divisor_n_reg_17_ ( .D(U17_Z_17), .CK(clock), .RN(n1206), .Q(
        U14_DATA1_17), .QN(n1125) );
  DFFR_X1 pipe2_divisor_n_reg_16_ ( .D(U17_Z_16), .CK(clock), .RN(n1198), .Q(
        U14_DATA1_16), .QN(n1162) );
  DFFR_X1 pipe2_divisor_n_reg_15_ ( .D(U17_Z_15), .CK(clock), .RN(n1200), .Q(
        U14_DATA1_15), .QN(n1121) );
  DFFR_X1 pipe2_divisor_n_reg_14_ ( .D(U17_Z_14), .CK(clock), .RN(n1201), .Q(
        U14_DATA1_14), .QN(n1117) );
  DFFR_X1 pipe2_divisor_n_reg_13_ ( .D(U17_Z_13), .CK(clock), .RN(n1201), .Q(
        U14_DATA1_13), .QN(n1113) );
  DFFR_X1 pipe2_divisor_n_reg_12_ ( .D(U17_Z_12), .CK(clock), .RN(n1203), .Q(
        U14_DATA1_12), .QN(n1159) );
  DFFR_X1 pipe2_divisor_n_reg_11_ ( .D(U17_Z_11), .CK(clock), .RN(n1204), .Q(
        U14_DATA1_11), .QN(n1109) );
  DFFR_X1 pipe2_divisor_n_reg_10_ ( .D(U17_Z_10), .CK(clock), .RN(n1205), .Q(
        U14_DATA1_10), .QN(n1155) );
  DFFR_X1 pipe2_divisor_n_reg_9_ ( .D(U17_Z_9), .CK(clock), .RN(n1207), .Q(
        U14_DATA1_9), .QN(n1105) );
  DFFR_X1 pipe2_divisor_n_reg_8_ ( .D(U17_Z_8), .CK(clock), .RN(n1208), .Q(
        U14_DATA1_8), .QN(n1151) );
  DFFR_X1 pipe2_divisor_n_reg_7_ ( .D(U17_Z_7), .CK(clock), .RN(n1185), .Q(
        U14_DATA1_7), .QN(n1101) );
  DFFR_X1 pipe2_divisor_n_reg_6_ ( .D(U17_Z_6), .CK(clock), .RN(n1188), .Q(
        U14_DATA1_6), .QN(n1097) );
  DFFR_X1 pipe2_divisor_n_reg_5_ ( .D(U17_Z_5), .CK(clock), .RN(n1190), .Q(
        U14_DATA1_5), .QN(n1093) );
  DFFR_X1 pipe2_divisor_n_reg_4_ ( .D(U17_Z_4), .CK(clock), .RN(n1194), .Q(
        U14_DATA1_4), .QN(n1147) );
  DFFR_X1 pipe2_divisor_n_reg_3_ ( .D(U17_Z_3), .CK(clock), .RN(n1199), .Q(
        U14_DATA1_3), .QN(n1089) );
  DFFR_X1 pipe2_divisor_n_reg_2_ ( .D(U17_Z_2), .CK(clock), .RN(n1202), .Q(
        U14_DATA1_2), .QN(n1143) );
  DFFR_X1 pipe2_divisor_n_reg_1_ ( .D(U17_Z_1), .CK(clock), .RN(n1198), .Q(
        U14_DATA1_1), .QN(n1085) );
  DFFR_X1 pipe2_divisor_n_reg_0_ ( .D(U17_Z_0), .CK(clock), .RN(n1204), .Q(
        U14_DATA1_0), .QN(n1138) );
  DFFR_X1 pipe2_result_reg_26_ ( .D(U18_Z_26), .CK(clock), .RN(n1199), .Q(n675) );
  DFFR_X1 pipe2_result_reg_25_ ( .D(U18_Z_25), .CK(clock), .RN(n1200), .Q(n674) );
  DFFR_X1 pipe2_result_reg_24_ ( .D(U18_Z_24), .CK(clock), .RN(n1195), .Q(n673) );
  DFFR_X1 pipe2_result_reg_23_ ( .D(U18_Z_23), .CK(clock), .RN(n1192), .Q(n672) );
  DFFR_X1 pipe2_result_reg_22_ ( .D(U18_Z_22), .CK(clock), .RN(n1204), .Q(n671) );
  DFFR_X1 pipe2_result_reg_21_ ( .D(U18_Z_21), .CK(clock), .RN(n1198), .Q(n670) );
  DFFR_X1 pipe2_result_reg_20_ ( .D(U18_Z_20), .CK(clock), .RN(n1200), .Q(n669) );
  DFFR_X1 pipe2_result_reg_19_ ( .D(U18_Z_19), .CK(clock), .RN(n1201), .Q(n668) );
  DFFR_X1 pipe2_result_reg_18_ ( .D(U18_Z_18), .CK(clock), .RN(n1203), .Q(n667) );
  DFFR_X1 pipe2_result_reg_17_ ( .D(U18_Z_17), .CK(clock), .RN(n1204), .Q(n666) );
  DFFR_X1 pipe2_result_reg_16_ ( .D(U18_Z_16), .CK(clock), .RN(n1205), .Q(n665) );
  DFFR_X1 pipe2_result_reg_15_ ( .D(U18_Z_15), .CK(clock), .RN(n1207), .Q(n664) );
  DFFR_X1 pipe2_result_reg_14_ ( .D(U18_Z_14), .CK(clock), .RN(n1208), .Q(n663) );
  DFFR_X1 pipe2_result_reg_13_ ( .D(U18_Z_13), .CK(clock), .RN(n1185), .Q(n662) );
  DFFR_X1 pipe2_result_reg_12_ ( .D(U18_Z_12), .CK(clock), .RN(n1188), .Q(n661) );
  DFFR_X1 pipe2_result_reg_11_ ( .D(U18_Z_11), .CK(clock), .RN(n1190), .Q(n660) );
  DFFR_X1 pipe2_result_reg_10_ ( .D(U18_Z_10), .CK(clock), .RN(n1194), .Q(n659) );
  DFFR_X1 pipe2_result_reg_9_ ( .D(U18_Z_9), .CK(clock), .RN(n1204), .Q(n658)
         );
  DFFR_X1 pipe2_result_reg_8_ ( .D(U18_Z_8), .CK(clock), .RN(n1205), .Q(n657)
         );
  DFFR_X1 pipe2_result_reg_7_ ( .D(U18_Z_7), .CK(clock), .RN(n1207), .Q(n656)
         );
  DFFR_X1 pipe2_result_reg_1_ ( .D(U18_Z_1), .CK(clock), .RN(n1208), .Q(n650)
         );
  DFFR_X1 pipe3_divisor_n_reg_19_ ( .D(U14_Z_19), .CK(clock), .RN(n1185), .Q(
        U11_DATA1_19) );
  DFFR_X1 pipe3_divisor_n_reg_18_ ( .D(U14_Z_18), .CK(clock), .RN(n1188), .Q(
        U11_DATA1_18), .QN(n1167) );
  DFFR_X1 pipe3_divisor_n_reg_17_ ( .D(U14_Z_17), .CK(clock), .RN(n1199), .Q(
        U11_DATA1_17), .QN(n1126) );
  DFFR_X1 pipe3_divisor_n_reg_16_ ( .D(U14_Z_16), .CK(clock), .RN(n1202), .Q(
        U11_DATA1_16), .QN(n1163) );
  DFFR_X1 pipe3_divisor_n_reg_15_ ( .D(U14_Z_15), .CK(clock), .RN(n1206), .Q(
        U11_DATA1_15), .QN(n1122) );
  DFFR_X1 pipe3_divisor_n_reg_14_ ( .D(U14_Z_14), .CK(clock), .RN(n1198), .Q(
        U11_DATA1_14), .QN(n1118) );
  DFFR_X1 pipe3_divisor_n_reg_13_ ( .D(U14_Z_13), .CK(clock), .RN(n1200), .Q(
        U11_DATA1_13), .QN(n1114) );
  DFFR_X1 pipe3_divisor_n_reg_12_ ( .D(U14_Z_12), .CK(clock), .RN(n1201), .Q(
        U11_DATA1_12), .QN(n1160) );
  DFFR_X1 pipe3_divisor_n_reg_11_ ( .D(U14_Z_11), .CK(clock), .RN(n1203), .Q(
        U11_DATA1_11), .QN(n1110) );
  DFFR_X1 pipe3_divisor_n_reg_10_ ( .D(U14_Z_10), .CK(clock), .RN(n1204), .Q(
        U11_DATA1_10), .QN(n1156) );
  DFFR_X1 pipe3_divisor_n_reg_9_ ( .D(U14_Z_9), .CK(clock), .RN(n1205), .Q(
        U11_DATA1_9), .QN(n1106) );
  DFFR_X1 pipe3_divisor_n_reg_8_ ( .D(U14_Z_8), .CK(clock), .RN(n1207), .Q(
        U11_DATA1_8), .QN(n1152) );
  DFFR_X1 pipe3_divisor_n_reg_7_ ( .D(U14_Z_7), .CK(clock), .RN(n1208), .Q(
        U11_DATA1_7), .QN(n1102) );
  DFFR_X1 pipe3_divisor_n_reg_6_ ( .D(U14_Z_6), .CK(clock), .RN(n1185), .Q(
        U11_DATA1_6), .QN(n1098) );
  DFFR_X1 pipe3_divisor_n_reg_5_ ( .D(U14_Z_5), .CK(clock), .RN(n1190), .Q(
        U11_DATA1_5), .QN(n1094) );
  DFFR_X1 pipe3_divisor_n_reg_4_ ( .D(U14_Z_4), .CK(clock), .RN(n1194), .Q(
        U11_DATA1_4), .QN(n1148) );
  DFFR_X1 pipe3_divisor_n_reg_3_ ( .D(U14_Z_3), .CK(clock), .RN(n1199), .Q(
        U11_DATA1_3), .QN(n1090) );
  DFFR_X1 pipe3_divisor_n_reg_2_ ( .D(U14_Z_2), .CK(clock), .RN(n1202), .Q(
        U11_DATA1_2), .QN(n1144) );
  DFFR_X1 pipe3_divisor_n_reg_1_ ( .D(U14_Z_1), .CK(clock), .RN(n1206), .Q(
        U11_DATA1_1), .QN(n1086) );
  DFFR_X1 pipe3_divisor_n_reg_0_ ( .D(U14_Z_0), .CK(clock), .RN(n1198), .Q(
        U11_DATA1_0), .QN(n1139) );
  DFFR_X1 pipe3_result_reg_26_ ( .D(U15_Z_26), .CK(clock), .RN(n1203), .Q(n542) );
  DFFR_X1 pipe3_result_reg_25_ ( .D(U15_Z_25), .CK(clock), .RN(n1204), .Q(n541) );
  DFFR_X1 pipe3_result_reg_24_ ( .D(U15_Z_24), .CK(clock), .RN(n1205), .Q(n540) );
  DFFR_X1 pipe3_result_reg_23_ ( .D(U15_Z_23), .CK(clock), .RN(n1207), .Q(n539) );
  DFFR_X1 pipe3_result_reg_22_ ( .D(U15_Z_22), .CK(clock), .RN(n1208), .Q(n538) );
  DFFR_X1 pipe3_result_reg_21_ ( .D(U15_Z_21), .CK(clock), .RN(n1185), .Q(n537) );
  DFFR_X1 pipe3_result_reg_20_ ( .D(U15_Z_20), .CK(clock), .RN(n1188), .Q(n536) );
  DFFR_X1 pipe3_result_reg_19_ ( .D(U15_Z_19), .CK(clock), .RN(n1190), .Q(n535) );
  DFFR_X1 pipe3_result_reg_18_ ( .D(U15_Z_18), .CK(clock), .RN(n1194), .Q(n534) );
  DFFR_X1 pipe3_result_reg_17_ ( .D(U15_Z_17), .CK(clock), .RN(n1199), .Q(n533) );
  DFFR_X1 pipe3_result_reg_16_ ( .D(U15_Z_16), .CK(clock), .RN(n1202), .Q(n532) );
  DFFR_X1 pipe3_result_reg_15_ ( .D(U15_Z_15), .CK(clock), .RN(n1206), .Q(n531) );
  DFFR_X1 pipe3_result_reg_14_ ( .D(U15_Z_14), .CK(clock), .RN(n1189), .Q(n530) );
  DFFR_X1 pipe3_result_reg_13_ ( .D(U15_Z_13), .CK(clock), .RN(n1189), .Q(n529) );
  DFFR_X1 pipe3_result_reg_12_ ( .D(U15_Z_12), .CK(clock), .RN(n1189), .Q(n528) );
  DFFR_X1 pipe3_result_reg_11_ ( .D(U15_Z_11), .CK(clock), .RN(n1189), .Q(n527) );
  DFFR_X1 pipe3_result_reg_10_ ( .D(U15_Z_10), .CK(clock), .RN(n1189), .Q(n526) );
  DFFR_X1 pipe3_result_reg_9_ ( .D(U15_Z_9), .CK(clock), .RN(n1189), .Q(n525)
         );
  DFFR_X1 pipe3_result_reg_8_ ( .D(U15_Z_8), .CK(clock), .RN(n1189), .Q(n524)
         );
  DFFR_X1 pipe3_result_reg_7_ ( .D(U15_Z_7), .CK(clock), .RN(n1189), .Q(n523)
         );
  DFFR_X1 pipe3_result_reg_1_ ( .D(U15_Z_1), .CK(clock), .RN(n1194), .Q(n517)
         );
  DFFR_X1 pipe4_divisor_n_reg_19_ ( .D(U11_Z_19), .CK(clock), .RN(n1199), .Q(
        U8_DATA1_19) );
  DFFR_X1 pipe4_divisor_n_reg_18_ ( .D(U11_Z_18), .CK(clock), .RN(n1202), .Q(
        U8_DATA1_18), .QN(n1168) );
  DFFR_X1 pipe4_divisor_n_reg_17_ ( .D(U11_Z_17), .CK(clock), .RN(n1206), .Q(
        U8_DATA1_17) );
  DFFR_X1 pipe4_divisor_n_reg_16_ ( .D(U11_Z_16), .CK(clock), .RN(n1198), .Q(
        U8_DATA1_16), .QN(n1164) );
  DFFR_X1 pipe4_divisor_n_reg_15_ ( .D(U11_Z_15), .CK(clock), .RN(n1200), .Q(
        U8_DATA1_15), .QN(n1123) );
  DFFR_X1 pipe4_divisor_n_reg_14_ ( .D(U11_Z_14), .CK(clock), .RN(n1201), .Q(
        U8_DATA1_14), .QN(n1119) );
  DFFR_X1 pipe4_divisor_n_reg_13_ ( .D(U11_Z_13), .CK(clock), .RN(n1203), .Q(
        U8_DATA1_13), .QN(n1115) );
  DFFR_X1 pipe4_divisor_n_reg_12_ ( .D(U11_Z_12), .CK(clock), .RN(n1204), .Q(
        U8_DATA1_12), .QN(n1161) );
  DFFR_X1 pipe4_divisor_n_reg_11_ ( .D(U11_Z_11), .CK(clock), .RN(n1205), .Q(
        U8_DATA1_11), .QN(n1111) );
  DFFR_X1 pipe4_divisor_n_reg_10_ ( .D(U11_Z_10), .CK(clock), .RN(n1189), .Q(
        U8_DATA1_10), .QN(n1157) );
  DFFR_X1 pipe4_divisor_n_reg_9_ ( .D(U11_Z_9), .CK(clock), .RN(n1189), .Q(
        U8_DATA1_9), .QN(n1107) );
  DFFR_X1 pipe4_divisor_n_reg_8_ ( .D(U11_Z_8), .CK(clock), .RN(n1189), .Q(
        U8_DATA1_8), .QN(n1153) );
  DFFR_X1 pipe4_divisor_n_reg_7_ ( .D(U11_Z_7), .CK(clock), .RN(n1189), .Q(
        U8_DATA1_7), .QN(n1103) );
  DFFR_X1 pipe4_divisor_n_reg_6_ ( .D(U11_Z_6), .CK(clock), .RN(n1189), .Q(
        U8_DATA1_6), .QN(n1099) );
  DFFR_X1 pipe4_divisor_n_reg_5_ ( .D(U11_Z_5), .CK(clock), .RN(n1197), .Q(
        U8_DATA1_5), .QN(n1095) );
  DFFR_X1 pipe4_divisor_n_reg_4_ ( .D(U11_Z_4), .CK(clock), .RN(n1209), .Q(
        U8_DATA1_4), .QN(n1149) );
  DFFR_X1 pipe4_divisor_n_reg_3_ ( .D(U11_Z_3), .CK(clock), .RN(n1189), .Q(
        U8_DATA1_3), .QN(n1091) );
  DFFR_X1 pipe4_divisor_n_reg_2_ ( .D(U11_Z_2), .CK(clock), .RN(n1191), .Q(
        U8_DATA1_2), .QN(n1145) );
  DFFR_X1 pipe4_divisor_n_reg_1_ ( .D(U11_Z_1), .CK(clock), .RN(n1186), .Q(
        U8_DATA1_1), .QN(n1087) );
  DFFR_X1 pipe4_divisor_n_reg_0_ ( .D(U11_Z_0), .CK(clock), .RN(n1187), .Q(
        U8_DATA1_0), .QN(n1140) );
  DFFR_X1 pipe4_result_reg_26_ ( .D(U12_Z_26), .CK(clock), .RN(n1193), .Q(n407) );
  DFFR_X1 pipe4_result_reg_25_ ( .D(U12_Z_25), .CK(clock), .RN(n1195), .Q(n406) );
  DFFR_X1 pipe4_result_reg_24_ ( .D(U12_Z_24), .CK(clock), .RN(n1196), .Q(n405) );
  DFFR_X1 pipe4_result_reg_23_ ( .D(U12_Z_23), .CK(clock), .RN(n1191), .Q(n404) );
  DFFR_X1 pipe4_result_reg_22_ ( .D(U12_Z_22), .CK(clock), .RN(n1186), .Q(n403) );
  DFFR_X1 pipe4_result_reg_21_ ( .D(U12_Z_21), .CK(clock), .RN(n1187), .Q(n402) );
  DFFR_X1 pipe4_result_reg_20_ ( .D(U12_Z_20), .CK(clock), .RN(n1200), .Q(n401) );
  DFFR_X1 pipe4_result_reg_19_ ( .D(U12_Z_19), .CK(clock), .RN(n1201), .Q(n400) );
  DFFR_X1 pipe4_result_reg_18_ ( .D(U12_Z_18), .CK(clock), .RN(n1203), .Q(n399) );
  DFFR_X1 pipe4_result_reg_17_ ( .D(U12_Z_17), .CK(clock), .RN(n1204), .Q(n398) );
  DFFR_X1 pipe4_result_reg_16_ ( .D(U12_Z_16), .CK(clock), .RN(n1205), .Q(n397) );
  DFFR_X1 pipe4_result_reg_15_ ( .D(U12_Z_15), .CK(clock), .RN(n1207), .Q(n396) );
  DFFR_X1 pipe4_result_reg_14_ ( .D(U12_Z_14), .CK(clock), .RN(n1208), .Q(n395) );
  DFFR_X1 pipe4_result_reg_13_ ( .D(U12_Z_13), .CK(clock), .RN(n1185), .Q(n394) );
  DFFR_X1 pipe4_result_reg_12_ ( .D(U12_Z_12), .CK(clock), .RN(n1188), .Q(n393) );
  DFFR_X1 pipe4_result_reg_11_ ( .D(U12_Z_11), .CK(clock), .RN(n1190), .Q(n392) );
  DFFR_X1 pipe4_result_reg_10_ ( .D(U12_Z_10), .CK(clock), .RN(n1194), .Q(n391) );
  DFFR_X1 pipe4_result_reg_9_ ( .D(U12_Z_9), .CK(clock), .RN(n1199), .Q(n390)
         );
  DFFR_X1 pipe4_result_reg_8_ ( .D(U12_Z_8), .CK(clock), .RN(n1207), .Q(n389)
         );
  DFFR_X1 pipe4_result_reg_7_ ( .D(U12_Z_7), .CK(clock), .RN(n1208), .Q(n388)
         );
  DFFR_X1 pipe4_result_reg_1_ ( .D(U12_Z_1), .CK(clock), .RN(n1185), .Q(n382)
         );
  DFFR_X1 pipe5_divisor_n_reg_19_ ( .D(U8_Z_19), .CK(clock), .RN(n1188), .Q(
        U5_DATA1_19) );
  DFFR_X1 pipe5_divisor_n_reg_18_ ( .D(U8_Z_18), .CK(clock), .RN(n1190), .Q(
        U5_DATA1_18), .QN(n1169) );
  DFFR_X1 pipe5_divisor_n_reg_16_ ( .D(U8_Z_16), .CK(clock), .RN(n1205), .Q(
        U5_DATA1_16), .QN(n1170) );
  DFFR_X1 pipe5_divisor_n_reg_15_ ( .D(U8_Z_15), .CK(clock), .RN(n1207), .Q(
        U5_DATA1_15), .QN(n1127) );
  DFFR_X1 pipe5_divisor_n_reg_14_ ( .D(U8_Z_14), .CK(clock), .RN(n1208), .Q(
        U5_DATA1_14), .QN(n1128) );
  DFFR_X1 pipe5_divisor_n_reg_13_ ( .D(U8_Z_13), .CK(clock), .RN(n1185), .Q(
        U5_DATA1_13), .QN(n1129) );
  DFFR_X1 pipe5_divisor_n_reg_12_ ( .D(U8_Z_12), .CK(clock), .RN(n1188), .Q(
        U5_DATA1_12), .QN(n1171) );
  DFFR_X1 pipe5_divisor_n_reg_11_ ( .D(U8_Z_11), .CK(clock), .RN(n1190), .Q(
        U5_DATA1_11), .QN(n1130) );
  DFFR_X1 pipe5_divisor_n_reg_10_ ( .D(U8_Z_10), .CK(clock), .RN(n1194), .Q(
        U5_DATA1_10), .QN(n1172) );
  DFFR_X1 pipe5_divisor_n_reg_9_ ( .D(U8_Z_9), .CK(clock), .RN(n1199), .Q(
        U5_DATA1_9), .QN(n1131) );
  DFFR_X1 pipe5_divisor_n_reg_8_ ( .D(U8_Z_8), .CK(clock), .RN(n1202), .Q(
        U5_DATA1_8), .QN(n1173) );
  DFFR_X1 pipe5_divisor_n_reg_7_ ( .D(U8_Z_7), .CK(clock), .RN(n1206), .Q(
        U5_DATA1_7), .QN(n1132) );
  DFFR_X1 pipe5_divisor_n_reg_6_ ( .D(U8_Z_6), .CK(clock), .RN(n1198), .Q(
        U5_DATA1_6), .QN(n1133) );
  DFFR_X1 pipe5_divisor_n_reg_5_ ( .D(U8_Z_5), .CK(clock), .RN(n1200), .Q(
        U5_DATA1_5), .QN(n1134) );
  DFFR_X1 pipe5_divisor_n_reg_4_ ( .D(U8_Z_4), .CK(clock), .RN(n1188), .Q(
        U5_DATA1_4), .QN(n1174) );
  DFFR_X1 pipe5_divisor_n_reg_3_ ( .D(U8_Z_3), .CK(clock), .RN(n1189), .Q(
        U5_DATA1_3), .QN(n1135) );
  DFFR_X1 pipe5_divisor_n_reg_2_ ( .D(U8_Z_2), .CK(clock), .RN(n1202), .Q(
        U5_DATA1_2), .QN(n1175) );
  DFFR_X1 pipe5_divisor_n_reg_1_ ( .D(U8_Z_1), .CK(clock), .RN(n1201), .Q(
        U5_DATA1_1), .QN(n1136) );
  DFFR_X1 pipe5_divisor_n_reg_0_ ( .D(U8_Z_0), .CK(clock), .RN(n1202), .Q(
        U5_DATA1_0), .QN(n1141) );
  DFFR_X1 pipe5_result_reg_26_ ( .D(U9_Z_26), .CK(clock), .RN(n1206), .Q(n270)
         );
  DFFR_X1 pipe5_result_reg_25_ ( .D(U9_Z_25), .CK(clock), .RN(n1201), .Q(n269)
         );
  DFFR_X1 pipe5_result_reg_24_ ( .D(U9_Z_24), .CK(clock), .RN(n1192), .Q(n268)
         );
  DFFR_X1 pipe5_result_reg_23_ ( .D(U9_Z_23), .CK(clock), .RN(n1200), .Q(n267)
         );
  DFFR_X1 pipe5_result_reg_22_ ( .D(U9_Z_22), .CK(clock), .RN(n1188), .Q(n266)
         );
  DFFR_X1 pipe5_result_reg_21_ ( .D(U9_Z_21), .CK(clock), .RN(n1204), .Q(n265)
         );
  DFFR_X1 pipe5_result_reg_20_ ( .D(U9_Z_20), .CK(clock), .RN(n1189), .Q(n264)
         );
  DFFR_X1 pipe5_result_reg_19_ ( .D(U9_Z_19), .CK(clock), .RN(n1194), .Q(n263)
         );
  DFFR_X1 pipe5_result_reg_18_ ( .D(U9_Z_18), .CK(clock), .RN(n1200), .Q(n262)
         );
  DFFR_X1 pipe5_result_reg_17_ ( .D(U9_Z_17), .CK(clock), .RN(n1201), .Q(n261)
         );
  DFFR_X1 pipe5_result_reg_16_ ( .D(U9_Z_16), .CK(clock), .RN(n1206), .Q(n260)
         );
  DFFR_X1 pipe5_result_reg_15_ ( .D(U9_Z_15), .CK(clock), .RN(n1203), .Q(n259)
         );
  DFFR_X1 pipe5_result_reg_14_ ( .D(U9_Z_14), .CK(clock), .RN(n1194), .Q(n258)
         );
  DFFR_X1 pipe5_result_reg_13_ ( .D(U9_Z_13), .CK(clock), .RN(n1201), .Q(n257)
         );
  DFFR_X1 pipe5_result_reg_12_ ( .D(U9_Z_12), .CK(clock), .RN(n1196), .Q(n256)
         );
  DFFR_X1 pipe5_result_reg_11_ ( .D(U9_Z_11), .CK(clock), .RN(n1193), .Q(n255)
         );
  DFFR_X1 pipe5_result_reg_10_ ( .D(U9_Z_10), .CK(clock), .RN(n1199), .Q(n254)
         );
  DFFR_X1 pipe5_result_reg_9_ ( .D(U9_Z_9), .CK(clock), .RN(n1203), .Q(n253)
         );
  DFFR_X1 pipe5_result_reg_8_ ( .D(U9_Z_8), .CK(clock), .RN(n1206), .Q(n252)
         );
  DFFR_X1 pipe5_result_reg_7_ ( .D(U9_Z_7), .CK(clock), .RN(n1190), .Q(n251)
         );
  DFFR_X1 pipe5_result_reg_1_ ( .D(U9_Z_1), .CK(clock), .RN(n1198), .Q(n245)
         );
  DFFR_X1 pipe6_result_reg_1_ ( .D(U6_Z_1), .CK(clock), .RN(n1203), .Q(n106)
         );
  INV_X4 U23 ( .A(divisor[19]), .ZN(n21) );
  AND2_X1 U46 ( .A1(U9_DATA1_6), .A2(n355), .ZN(U9_Z_6) );
  AND2_X1 U47 ( .A1(U9_DATA1_5), .A2(n355), .ZN(U9_Z_5) );
  AND2_X1 U48 ( .A1(U9_DATA1_4), .A2(n355), .ZN(U9_Z_4) );
  AND2_X1 U49 ( .A1(U9_DATA1_3), .A2(n355), .ZN(U9_Z_3) );
  AND2_X1 U58 ( .A1(U9_DATA1_2), .A2(n355), .ZN(U9_Z_2) );
  AND2_X1 U69 ( .A1(U9_DATA1_1), .A2(n355), .ZN(U9_Z_1) );
  AND2_X1 U79 ( .A1(U8_DATA1_19), .A2(n355), .ZN(U8_Z_19) );
  AND2_X1 U91 ( .A1(U7_DATA1_5), .A2(n355), .ZN(U7_Z_5) );
  AND2_X1 U92 ( .A1(U7_DATA1_4), .A2(n355), .ZN(U7_Z_4) );
  AND2_X1 U93 ( .A1(U7_DATA1_3), .A2(n355), .ZN(U7_Z_3) );
  AND2_X1 U94 ( .A1(U7_DATA1_2), .A2(n355), .ZN(U7_Z_2) );
  AND2_X1 U99 ( .A1(U6_DATA1_7), .A2(n217), .ZN(U6_Z_7) );
  AND2_X1 U100 ( .A1(U6_DATA1_6), .A2(n217), .ZN(U6_Z_6) );
  AND2_X1 U101 ( .A1(U6_DATA1_5), .A2(n217), .ZN(U6_Z_5) );
  AND2_X1 U102 ( .A1(U6_DATA1_4), .A2(n217), .ZN(U6_Z_4) );
  AND2_X1 U103 ( .A1(U6_DATA1_3), .A2(n217), .ZN(U6_Z_3) );
  AND2_X1 U112 ( .A1(U6_DATA1_2), .A2(n217), .ZN(U6_Z_2) );
  AND2_X1 U123 ( .A1(U6_DATA1_1), .A2(n217), .ZN(U6_Z_1) );
  AND2_X1 U133 ( .A1(U5_DATA1_19), .A2(n217), .ZN(U5_Z_19) );
  AND2_X1 U145 ( .A1(U4_DATA1_6), .A2(n217), .ZN(U4_Z_6) );
  AND2_X1 U146 ( .A1(U4_DATA1_5), .A2(n217), .ZN(U4_Z_5) );
  AND2_X1 U147 ( .A1(U4_DATA1_4), .A2(n217), .ZN(U4_Z_4) );
  AND2_X1 U148 ( .A1(U4_DATA1_3), .A2(n217), .ZN(U4_Z_3) );
  AND2_X1 U149 ( .A1(U4_DATA1_2), .A2(n217), .ZN(U4_Z_2) );
  AND2_X1 U155 ( .A1(U24_DATA1_6), .A2(start), .ZN(U24_Z_6) );
  AND2_X1 U156 ( .A1(U24_DATA1_5), .A2(start), .ZN(U24_Z_5) );
  AND2_X1 U157 ( .A1(U24_DATA1_4), .A2(start), .ZN(U24_Z_4) );
  AND2_X1 U158 ( .A1(U24_DATA1_3), .A2(start), .ZN(U24_Z_3) );
  AND2_X1 U167 ( .A1(U24_DATA1_2), .A2(start), .ZN(U24_Z_2) );
  AND2_X1 U178 ( .A1(U24_DATA1_1), .A2(n1183), .ZN(U24_Z_1) );
  AND2_X1 U184 ( .A1(U21_DATA1_6), .A2(n887), .ZN(U21_Z_6) );
  AND2_X1 U185 ( .A1(U21_DATA1_5), .A2(n887), .ZN(U21_Z_5) );
  AND2_X1 U186 ( .A1(U21_DATA1_4), .A2(n887), .ZN(U21_Z_4) );
  AND2_X1 U187 ( .A1(U21_DATA1_3), .A2(n887), .ZN(U21_Z_3) );
  AND2_X1 U196 ( .A1(U21_DATA1_2), .A2(n887), .ZN(U21_Z_2) );
  AND2_X1 U207 ( .A1(U21_DATA1_1), .A2(n887), .ZN(U21_Z_1) );
  AND2_X1 U217 ( .A1(U20_DATA1_19), .A2(n887), .ZN(U20_Z_19) );
  AND2_X1 U234 ( .A1(U18_DATA1_6), .A2(n1068), .ZN(U18_Z_6) );
  AND2_X1 U235 ( .A1(U18_DATA1_5), .A2(n1068), .ZN(U18_Z_5) );
  AND2_X1 U236 ( .A1(U18_DATA1_4), .A2(n1068), .ZN(U18_Z_4) );
  AND2_X1 U237 ( .A1(U18_DATA1_3), .A2(n1068), .ZN(U18_Z_3) );
  AND2_X1 U246 ( .A1(U18_DATA1_2), .A2(n1068), .ZN(U18_Z_2) );
  AND2_X1 U257 ( .A1(U18_DATA1_1), .A2(n1068), .ZN(U18_Z_1) );
  AND2_X1 U267 ( .A1(U17_DATA1_19), .A2(n1068), .ZN(U17_Z_19) );
  AND2_X1 U279 ( .A1(U16_DATA1_2), .A2(n1068), .ZN(U16_Z_2) );
  AND2_X1 U285 ( .A1(U15_DATA1_6), .A2(n625), .ZN(U15_Z_6) );
  AND2_X1 U286 ( .A1(U15_DATA1_5), .A2(n625), .ZN(U15_Z_5) );
  AND2_X1 U287 ( .A1(U15_DATA1_4), .A2(n625), .ZN(U15_Z_4) );
  AND2_X1 U288 ( .A1(U15_DATA1_3), .A2(n625), .ZN(U15_Z_3) );
  AND2_X1 U297 ( .A1(U15_DATA1_2), .A2(n625), .ZN(U15_Z_2) );
  AND2_X1 U308 ( .A1(U15_DATA1_1), .A2(n625), .ZN(U15_Z_1) );
  AND2_X1 U318 ( .A1(U14_DATA1_19), .A2(n625), .ZN(U14_Z_19) );
  AND2_X1 U330 ( .A1(U13_DATA1_3), .A2(n625), .ZN(U13_Z_3) );
  AND2_X1 U331 ( .A1(U13_DATA1_2), .A2(n625), .ZN(U13_Z_2) );
  AND2_X1 U337 ( .A1(U12_DATA1_6), .A2(n491), .ZN(U12_Z_6) );
  AND2_X1 U338 ( .A1(U12_DATA1_5), .A2(n491), .ZN(U12_Z_5) );
  AND2_X1 U339 ( .A1(U12_DATA1_4), .A2(n491), .ZN(U12_Z_4) );
  AND2_X1 U340 ( .A1(U12_DATA1_3), .A2(n491), .ZN(U12_Z_3) );
  AND2_X1 U349 ( .A1(U12_DATA1_2), .A2(n491), .ZN(U12_Z_2) );
  AND2_X1 U360 ( .A1(U12_DATA1_1), .A2(n491), .ZN(U12_Z_1) );
  AND2_X1 U370 ( .A1(U11_DATA1_19), .A2(n491), .ZN(U11_Z_19) );
  AND2_X1 U382 ( .A1(U10_DATA1_4), .A2(n491), .ZN(U10_Z_4) );
  AND2_X1 U383 ( .A1(U10_DATA1_3), .A2(n491), .ZN(U10_Z_3) );
  AND2_X1 U384 ( .A1(U10_DATA1_2), .A2(n491), .ZN(U10_Z_2) );
  DFFR_X2 StartOut1_reg ( .D(n887), .CK(clock), .RN(n1193), .Q(n1068), .QN(
        n1063) );
  DFFR_X2 StartOut0_reg ( .D(start), .CK(clock), .RN(n1191), .Q(n887), .QN(
        n1182) );
  DFFR_X2 pipe6_divisor_n_reg_4_ ( .D(U5_Z_4), .CK(clock), .RN(n1186), .Q(
        n[89]) );
  DFFR_X2 pipe6_divisor_n_reg_2_ ( .D(U5_Z_2), .CK(clock), .RN(n1197), .Q(
        n[87]) );
  DFFR_X2 pipe6_divisor_n_reg_0_ ( .D(U5_Z_0), .CK(clock), .RN(n1195), .Q(
        n[85]) );
  DFFR_X2 pipe6_divisor_n_reg_3_ ( .D(U5_Z_3), .CK(clock), .RN(n1186), .Q(
        n[88]) );
  DFFR_X2 pipe6_divisor_n_reg_1_ ( .D(U5_Z_1), .CK(clock), .RN(n1187), .Q(
        n[86]) );
  DFFR_X2 pipe6_divisor_n_reg_18_ ( .D(U5_Z_18), .CK(clock), .RN(n1189), .Q(
        n[103]) );
  DFFR_X2 pipe6_divisor_n_reg_17_ ( .D(U5_Z_17), .CK(clock), .RN(n1191), .Q(
        n[102]) );
  DFFR_X2 pipe6_divisor_n_reg_16_ ( .D(U5_Z_16), .CK(clock), .RN(n1186), .Q(
        n[101]) );
  DFFR_X2 pipe6_divisor_n_reg_15_ ( .D(U5_Z_15), .CK(clock), .RN(n1187), .Q(
        n[100]) );
  DFFR_X2 pipe6_divisor_n_reg_14_ ( .D(U5_Z_14), .CK(clock), .RN(n1192), .Q(
        n[99]) );
  DFFR_X2 pipe6_divisor_n_reg_13_ ( .D(U5_Z_13), .CK(clock), .RN(n1193), .Q(
        n[98]) );
  DFFR_X2 pipe6_divisor_n_reg_12_ ( .D(U5_Z_12), .CK(clock), .RN(n1195), .Q(
        n[97]) );
  DFFR_X2 pipe6_divisor_n_reg_11_ ( .D(U5_Z_11), .CK(clock), .RN(n1209), .Q(
        n[96]) );
  DFFR_X2 pipe6_divisor_n_reg_10_ ( .D(U5_Z_10), .CK(clock), .RN(n1196), .Q(
        n[95]) );
  DFFR_X2 pipe6_divisor_n_reg_9_ ( .D(U5_Z_9), .CK(clock), .RN(n1197), .Q(
        n[94]) );
  DFFR_X2 pipe6_divisor_n_reg_8_ ( .D(U5_Z_8), .CK(clock), .RN(n1191), .Q(
        n[93]) );
  DFFR_X2 pipe6_divisor_n_reg_7_ ( .D(U5_Z_7), .CK(clock), .RN(n1192), .Q(
        n[92]) );
  DFFR_X2 pipe6_divisor_n_reg_6_ ( .D(U5_Z_6), .CK(clock), .RN(n1191), .Q(
        n[91]) );
  DFFR_X2 pipe6_divisor_n_reg_5_ ( .D(U5_Z_5), .CK(clock), .RN(reset_n), .Q(
        n[90]) );
  DFFR_X2 pipe1_result_reg_6_ ( .D(U21_Z_6), .CK(clock), .RN(n1189), .Q(n786)
         );
  DFFR_X2 pipe1_result_reg_5_ ( .D(U21_Z_5), .CK(clock), .RN(n1192), .Q(n785)
         );
  DFFR_X2 pipe1_result_reg_4_ ( .D(U21_Z_4), .CK(clock), .RN(n1193), .Q(n784)
         );
  DFFR_X2 pipe1_result_reg_3_ ( .D(U21_Z_3), .CK(clock), .RN(n1195), .Q(n783)
         );
  DFFR_X2 pipe1_result_reg_2_ ( .D(U21_Z_2), .CK(clock), .RN(n1196), .Q(n782)
         );
  DFFR_X2 pipe1_q_reg_7_ ( .D(U19_Z_1), .CK(clock), .RN(n1192), .Q(U16_DATA1_2) );
  DFFR_X2 pipe0_result_reg_6_ ( .D(U24_Z_6), .CK(clock), .RN(n1209), .Q(n915)
         );
  DFFR_X2 pipe0_result_reg_5_ ( .D(U24_Z_5), .CK(clock), .RN(n1189), .Q(n914)
         );
  DFFR_X2 pipe0_result_reg_4_ ( .D(U24_Z_4), .CK(clock), .RN(n1191), .Q(n913)
         );
  DFFR_X2 pipe0_result_reg_3_ ( .D(U24_Z_3), .CK(clock), .RN(n1186), .Q(n912)
         );
  DFFR_X2 pipe0_result_reg_2_ ( .D(U24_Z_2), .CK(clock), .RN(n1197), .Q(n911)
         );
  DFFR_X2 pipe0_result_reg_1_ ( .D(U24_Z_1), .CK(clock), .RN(n1209), .Q(n910)
         );
  DFFR_X2 StartOut_reg ( .D(n217), .CK(clock), .RN(n1196), .Q(StartOut) );
  DFFR_X2 StartOut5_reg ( .D(n355), .CK(clock), .RN(n1189), .Q(n217), .QN(
        n1066) );
  DFFR_X2 StartOut4_reg ( .D(n491), .CK(clock), .RN(n1209), .Q(n355), .QN(
        n1067) );
  DFFR_X2 StartOut3_reg ( .D(n625), .CK(clock), .RN(n1193), .Q(n491), .QN(
        n1065) );
  DFFR_X2 StartOut2_reg ( .D(n1068), .CK(clock), .RN(n1186), .Q(n625), .QN(
        n1064) );
  DFFR_X2 pipe6_result_reg_7_ ( .D(U6_Z_7), .CK(clock), .RN(n1191), .Q(n112)
         );
  DFFR_X2 pipe6_result_reg_6_ ( .D(U6_Z_6), .CK(clock), .RN(n1186), .Q(n111)
         );
  DFFR_X2 pipe6_result_reg_5_ ( .D(U6_Z_5), .CK(clock), .RN(n1187), .Q(n110)
         );
  DFFR_X2 pipe6_result_reg_4_ ( .D(U6_Z_4), .CK(clock), .RN(n1192), .Q(n109)
         );
  DFFR_X2 pipe6_result_reg_3_ ( .D(U6_Z_3), .CK(clock), .RN(n1193), .Q(n108)
         );
  DFFR_X2 pipe6_result_reg_2_ ( .D(U6_Z_2), .CK(clock), .RN(n1195), .Q(n107)
         );
  DFFR_X2 pipe6_q_reg_7_ ( .D(U4_Z_6), .CK(clock), .RN(n1197), .Q(q[7]) );
  DFFR_X2 pipe6_q_reg_6_ ( .D(U4_Z_5), .CK(clock), .RN(n1209), .Q(q[6]) );
  DFFR_X2 pipe6_q_reg_5_ ( .D(U4_Z_4), .CK(clock), .RN(n1189), .Q(q[5]) );
  DFFR_X2 pipe6_q_reg_4_ ( .D(U4_Z_3), .CK(clock), .RN(n1191), .Q(q[4]) );
  DFFR_X2 pipe6_q_reg_3_ ( .D(U4_Z_2), .CK(clock), .RN(n1209), .Q(q[3]) );
  DFFR_X2 pipe6_q_reg_2_ ( .D(U4_Z_1), .CK(clock), .RN(n1186), .Q(q[2]) );
  DFFR_X2 pipe6_divisor_n_reg_19_ ( .D(U5_Z_19), .CK(clock), .RN(n1196), .Q(
        n[104]) );
  DFFR_X2 pipe5_result_reg_6_ ( .D(U9_Z_6), .CK(clock), .RN(n1189), .Q(n250)
         );
  DFFR_X2 pipe5_result_reg_5_ ( .D(U9_Z_5), .CK(clock), .RN(n1189), .Q(n249)
         );
  DFFR_X2 pipe5_result_reg_4_ ( .D(U9_Z_4), .CK(clock), .RN(n1209), .Q(n248)
         );
  DFFR_X2 pipe5_result_reg_3_ ( .D(U9_Z_3), .CK(clock), .RN(n1197), .Q(n247)
         );
  DFFR_X2 pipe5_result_reg_2_ ( .D(U9_Z_2), .CK(clock), .RN(n1209), .Q(n246)
         );
  DFFR_X2 pipe5_q_reg_7_ ( .D(U7_Z_5), .CK(clock), .RN(n1187), .Q(U4_DATA1_6)
         );
  DFFR_X2 pipe5_q_reg_6_ ( .D(U7_Z_4), .CK(clock), .RN(n1197), .Q(U4_DATA1_5)
         );
  DFFR_X2 pipe5_q_reg_5_ ( .D(U7_Z_3), .CK(clock), .RN(n1191), .Q(U4_DATA1_4)
         );
  DFFR_X2 pipe5_q_reg_4_ ( .D(U7_Z_2), .CK(clock), .RN(n1191), .Q(U4_DATA1_3)
         );
  DFFR_X2 pipe5_q_reg_3_ ( .D(U7_Z_1), .CK(clock), .RN(n1189), .Q(U4_DATA1_2)
         );
  DFFR_X2 pipe4_result_reg_6_ ( .D(U12_Z_6), .CK(clock), .RN(n1192), .Q(n387)
         );
  DFFR_X2 pipe4_result_reg_5_ ( .D(U12_Z_5), .CK(clock), .RN(n1193), .Q(n386)
         );
  DFFR_X2 pipe4_result_reg_4_ ( .D(U12_Z_4), .CK(clock), .RN(n1195), .Q(n385)
         );
  DFFR_X2 pipe4_result_reg_3_ ( .D(U12_Z_3), .CK(clock), .RN(n1196), .Q(n384)
         );
  DFFR_X2 pipe4_result_reg_2_ ( .D(U12_Z_2), .CK(clock), .RN(n1197), .Q(n383)
         );
  DFFR_X2 pipe4_q_reg_7_ ( .D(U10_Z_4), .CK(clock), .RN(n1197), .Q(U7_DATA1_5)
         );
  DFFR_X2 pipe4_q_reg_6_ ( .D(U10_Z_3), .CK(clock), .RN(n1191), .Q(U7_DATA1_4)
         );
  DFFR_X2 pipe4_q_reg_5_ ( .D(U10_Z_2), .CK(clock), .RN(n1186), .Q(U7_DATA1_3)
         );
  DFFR_X2 pipe4_q_reg_4_ ( .D(U10_Z_1), .CK(clock), .RN(n1187), .Q(U7_DATA1_2)
         );
  DFFR_X2 pipe3_result_reg_6_ ( .D(U15_Z_6), .CK(clock), .RN(n1187), .Q(n522)
         );
  DFFR_X2 pipe3_result_reg_5_ ( .D(U15_Z_5), .CK(clock), .RN(n1192), .Q(n521)
         );
  DFFR_X2 pipe3_result_reg_4_ ( .D(U15_Z_4), .CK(clock), .RN(n1193), .Q(n520)
         );
  DFFR_X2 pipe3_result_reg_3_ ( .D(U15_Z_3), .CK(clock), .RN(n1195), .Q(n519)
         );
  DFFR_X2 pipe3_result_reg_2_ ( .D(U15_Z_2), .CK(clock), .RN(n1191), .Q(n518)
         );
  DFFR_X2 pipe3_q_reg_7_ ( .D(U13_Z_3), .CK(clock), .RN(n1195), .Q(U10_DATA1_4) );
  DFFR_X2 pipe3_q_reg_6_ ( .D(U13_Z_2), .CK(clock), .RN(n1196), .Q(U10_DATA1_3) );
  DFFR_X2 pipe3_q_reg_5_ ( .D(U13_Z_1), .CK(clock), .RN(n1197), .Q(U10_DATA1_2) );
  DFFR_X2 pipe2_result_reg_6_ ( .D(U18_Z_6), .CK(clock), .RN(n1186), .Q(n655)
         );
  DFFR_X2 pipe2_result_reg_5_ ( .D(U18_Z_5), .CK(clock), .RN(n1187), .Q(n654)
         );
  DFFR_X2 pipe2_result_reg_4_ ( .D(U18_Z_4), .CK(clock), .RN(n1192), .Q(n653)
         );
  DFFR_X2 pipe2_result_reg_3_ ( .D(U18_Z_3), .CK(clock), .RN(n1193), .Q(n652)
         );
  DFFR_X2 pipe2_result_reg_2_ ( .D(U18_Z_2), .CK(clock), .RN(n1195), .Q(n651)
         );
  DFFR_X2 pipe2_q_reg_7_ ( .D(U16_Z_2), .CK(clock), .RN(n1192), .Q(U13_DATA1_3) );
  DFFR_X2 pipe2_q_reg_6_ ( .D(U16_Z_1), .CK(clock), .RN(n1209), .Q(U13_DATA1_2) );
  DFFR_X2 pipe1_q_reg_6_ ( .D(U19_Z_0), .CK(clock), .RN(n1196), .Q(U16_DATA1_1) );
  DFFR_X2 pipe0_q_reg_7_ ( .D(U22_Z_0), .CK(clock), .RN(n1186), .Q(U19_DATA1_1) );
  DFFR_X2 pipe6_q_reg_1_ ( .D(U4_Z_0), .CK(clock), .RN(n1187), .Q(q[1]) );
  DFFR_X2 pipe5_q_reg_2_ ( .D(U7_Z_0), .CK(clock), .RN(n1209), .Q(U4_DATA1_1)
         );
  DFFR_X2 pipe4_q_reg_3_ ( .D(U10_Z_0), .CK(clock), .RN(n1193), .Q(U7_DATA1_1)
         );
  DFFR_X2 pipe3_q_reg_4_ ( .D(U13_Z_0), .CK(clock), .RN(n1209), .Q(U10_DATA1_1) );
  DFFR_X2 pipe2_q_reg_5_ ( .D(U16_Z_0), .CK(clock), .RN(n1196), .Q(U13_DATA1_1) );
  DFFR_X2 pipe2_divisor_n_reg_19_ ( .D(U17_Z_19), .CK(clock), .RN(n1189), .Q(
        U14_DATA1_19) );
  DFFR_X2 pipe1_divisor_n_reg_16_ ( .D(U20_Z_16), .CK(clock), .RN(n1186), .Q(
        U17_DATA1_16), .QN(n1214) );
  SDFFR_X1 pipe0_divisor_n_reg_19_ ( .D(start), .SI(1'b0), .SE(divisor[19]), 
        .CK(clock), .RN(reset_n), .Q(U20_DATA1_19) );
  DFFR_X2 pipe0_divisor_n_reg_1_ ( .D(n1180), .CK(clock), .RN(n1187), .Q(
        U20_DATA1_1), .QN(n1210) );
  DFFR_X2 pipe0_divisor_n_reg_3_ ( .D(n1179), .CK(clock), .RN(n1192), .Q(
        U20_DATA1_3), .QN(n1211) );
  DFFR_X2 pipe0_divisor_n_reg_9_ ( .D(n1178), .CK(clock), .RN(n1193), .Q(
        U20_DATA1_9), .QN(n1212) );
  DFFR_X2 pipe0_divisor_n_reg_11_ ( .D(n1177), .CK(clock), .RN(n1195), .Q(
        U20_DATA1_11), .QN(n1213) );
  SDFFR_X1 pipe5_divisor_n_reg_17_ ( .D(1'b0), .SI(U8_DATA1_17), .SE(n355), 
        .CK(clock), .RN(reset_n), .Q(U5_DATA1_17), .QN(n1215) );
  DFFR_X2 pipe1_result_reg_27_ ( .D(U21_Z_27), .CK(clock), .RN(n1197), .Q(n807) );
  DFFR_X2 pipe0_result_reg_27_ ( .D(U24_Z_27), .CK(clock), .RN(n1196), .Q(n936) );
  DFFR_X2 pipe6_result_reg_26_ ( .D(U6_Z_26), .CK(clock), .RN(n1192), .Q(n131)
         );
  DFFR_X2 pipe6_result_reg_25_ ( .D(U6_Z_25), .CK(clock), .RN(n1193), .Q(n130)
         );
  DFFR_X2 pipe6_result_reg_24_ ( .D(U6_Z_24), .CK(clock), .RN(n1195), .Q(n129)
         );
  DFFR_X2 pipe6_result_reg_23_ ( .D(U6_Z_23), .CK(clock), .RN(n1197), .Q(n128)
         );
  DFFR_X2 pipe6_result_reg_22_ ( .D(U6_Z_22), .CK(clock), .RN(n1189), .Q(n127)
         );
  DFFR_X2 pipe6_result_reg_21_ ( .D(U6_Z_21), .CK(clock), .RN(n1191), .Q(n126)
         );
  DFFR_X2 pipe6_result_reg_20_ ( .D(U6_Z_20), .CK(clock), .RN(n1209), .Q(n125)
         );
  DFFR_X2 pipe6_result_reg_19_ ( .D(U6_Z_19), .CK(clock), .RN(n1186), .Q(n124)
         );
  DFFR_X2 pipe6_result_reg_18_ ( .D(U6_Z_18), .CK(clock), .RN(n1187), .Q(n123)
         );
  DFFR_X2 pipe6_result_reg_17_ ( .D(U6_Z_17), .CK(clock), .RN(n1192), .Q(n122)
         );
  DFFR_X2 pipe6_result_reg_16_ ( .D(U6_Z_16), .CK(clock), .RN(n1193), .Q(n121)
         );
  DFFR_X2 pipe6_result_reg_15_ ( .D(U6_Z_15), .CK(clock), .RN(n1195), .Q(n120)
         );
  DFFR_X2 pipe6_result_reg_14_ ( .D(U6_Z_14), .CK(clock), .RN(n1196), .Q(n119)
         );
  DFFR_X2 pipe6_result_reg_13_ ( .D(U6_Z_13), .CK(clock), .RN(n1197), .Q(n118)
         );
  DFFR_X2 pipe6_result_reg_12_ ( .D(U6_Z_12), .CK(clock), .RN(n1189), .Q(n117)
         );
  DFFR_X2 pipe6_result_reg_11_ ( .D(U6_Z_11), .CK(clock), .RN(n1196), .Q(n116)
         );
  DFFR_X2 pipe6_result_reg_27_ ( .D(U6_Z_27), .CK(clock), .RN(n1196), .Q(n132)
         );
  DFFR_X2 pipe6_result_reg_10_ ( .D(U6_Z_10), .CK(clock), .RN(n1197), .Q(n115)
         );
  DFFR_X2 pipe6_result_reg_9_ ( .D(U6_Z_9), .CK(clock), .RN(n1209), .Q(n114)
         );
  DFFR_X2 pipe6_result_reg_8_ ( .D(U6_Z_8), .CK(clock), .RN(n1189), .Q(n113)
         );
  DFFR_X2 pipe5_result_reg_27_ ( .D(U9_Z_27), .CK(clock), .RN(n1187), .Q(n271)
         );
  DFFR_X2 pipe4_result_reg_27_ ( .D(U12_Z_27), .CK(clock), .RN(n1195), .Q(n408) );
  DFFR_X2 pipe3_result_reg_27_ ( .D(U15_Z_27), .CK(clock), .RN(n1189), .Q(n543) );
  DFFR_X2 pipe2_result_reg_27_ ( .D(U18_Z_27), .CK(clock), .RN(n1187), .Q(n676) );
  AND2_X1 U6 ( .A1(n1223), .A2(start), .ZN(n1177) );
  AND2_X1 U12 ( .A1(n1225), .A2(start), .ZN(n1178) );
  AND2_X1 U14 ( .A1(n1231), .A2(n1183), .ZN(n1179) );
  AND2_X1 U22 ( .A1(n1233), .A2(n1183), .ZN(n1180) );
  INV_X4 U25 ( .A(n1184), .ZN(n1183) );
  BUF_X4 U26 ( .A(reset_n), .Z(n1186) );
  BUF_X4 U27 ( .A(reset_n), .Z(n1187) );
  BUF_X4 U29 ( .A(reset_n), .Z(n1191) );
  BUF_X4 U30 ( .A(reset_n), .Z(n1192) );
  BUF_X4 U31 ( .A(reset_n), .Z(n1193) );
  BUF_X4 U32 ( .A(reset_n), .Z(n1195) );
  BUF_X4 U33 ( .A(reset_n), .Z(n1196) );
  BUF_X4 U34 ( .A(reset_n), .Z(n1197) );
  BUF_X4 U35 ( .A(reset_n), .Z(n1198) );
  BUF_X4 U36 ( .A(reset_n), .Z(n1200) );
  BUF_X4 U37 ( .A(reset_n), .Z(n1201) );
  BUF_X4 U38 ( .A(reset_n), .Z(n1203) );
  BUF_X4 U39 ( .A(reset_n), .Z(n1204) );
  BUF_X4 U40 ( .A(reset_n), .Z(n1205) );
  BUF_X4 U41 ( .A(reset_n), .Z(n1207) );
  BUF_X4 U42 ( .A(reset_n), .Z(n1208) );
  BUF_X4 U43 ( .A(reset_n), .Z(n1209) );
  BUF_X4 U44 ( .A(reset_n), .Z(n1185) );
  BUF_X4 U45 ( .A(reset_n), .Z(n1188) );
  BUF_X4 U50 ( .A(reset_n), .Z(n1190) );
  BUF_X4 U51 ( .A(reset_n), .Z(n1194) );
  BUF_X4 U52 ( .A(reset_n), .Z(n1199) );
  BUF_X4 U53 ( .A(reset_n), .Z(n1202) );
  BUF_X4 U54 ( .A(reset_n), .Z(n1206) );
  INV_X4 U55 ( .A(start), .ZN(n1184) );
  INV_X4 U64 ( .A(divisor[0]), .ZN(n1234) );
  NOR2_X2 U65 ( .A1(n1182), .A2(n1077), .ZN(U20_Z_0) );
  NOR2_X2 U66 ( .A1(n1063), .A2(n1137), .ZN(U17_Z_0) );
  NOR2_X2 U67 ( .A1(n1064), .A2(n1138), .ZN(U14_Z_0) );
  NOR2_X2 U68 ( .A1(n1065), .A2(n1139), .ZN(U11_Z_0) );
  NOR2_X2 U70 ( .A1(n1067), .A2(n1140), .ZN(U8_Z_0) );
  INV_X4 U71 ( .A(divisor[1]), .ZN(n1233) );
  NOR2_X2 U72 ( .A1(n1182), .A2(n1210), .ZN(U20_Z_1) );
  NOR2_X2 U73 ( .A1(n1063), .A2(n1084), .ZN(U17_Z_1) );
  NOR2_X2 U74 ( .A1(n1064), .A2(n1085), .ZN(U14_Z_1) );
  NOR2_X2 U75 ( .A1(n1065), .A2(n1086), .ZN(U11_Z_1) );
  NOR2_X2 U76 ( .A1(n1067), .A2(n1087), .ZN(U8_Z_1) );
  INV_X4 U77 ( .A(divisor[2]), .ZN(n1232) );
  NOR2_X2 U78 ( .A1(n1182), .A2(n1078), .ZN(U20_Z_2) );
  NOR2_X2 U80 ( .A1(n1063), .A2(n1142), .ZN(U17_Z_2) );
  NOR2_X2 U81 ( .A1(n1064), .A2(n1143), .ZN(U14_Z_2) );
  NOR2_X2 U82 ( .A1(n1065), .A2(n1144), .ZN(U11_Z_2) );
  NOR2_X2 U83 ( .A1(n1067), .A2(n1145), .ZN(U8_Z_2) );
  INV_X4 U84 ( .A(divisor[3]), .ZN(n1231) );
  NOR2_X2 U85 ( .A1(n1182), .A2(n1211), .ZN(U20_Z_3) );
  NOR2_X2 U86 ( .A1(n1063), .A2(n1088), .ZN(U17_Z_3) );
  NOR2_X2 U87 ( .A1(n1064), .A2(n1089), .ZN(U14_Z_3) );
  NOR2_X2 U88 ( .A1(n1065), .A2(n1090), .ZN(U11_Z_3) );
  NOR2_X2 U89 ( .A1(n1067), .A2(n1091), .ZN(U8_Z_3) );
  INV_X4 U90 ( .A(divisor[4]), .ZN(n1230) );
  NOR2_X2 U95 ( .A1(n1182), .A2(n1079), .ZN(U20_Z_4) );
  NOR2_X2 U96 ( .A1(n1063), .A2(n1146), .ZN(U17_Z_4) );
  NOR2_X2 U97 ( .A1(n1064), .A2(n1147), .ZN(U14_Z_4) );
  NOR2_X2 U98 ( .A1(n1065), .A2(n1148), .ZN(U11_Z_4) );
  NOR2_X2 U104 ( .A1(n1067), .A2(n1149), .ZN(U8_Z_4) );
  INV_X4 U105 ( .A(divisor[5]), .ZN(n1229) );
  NOR2_X2 U106 ( .A1(n1182), .A2(n1069), .ZN(U20_Z_5) );
  NOR2_X2 U107 ( .A1(n1063), .A2(n1092), .ZN(U17_Z_5) );
  NOR2_X2 U108 ( .A1(n1064), .A2(n1093), .ZN(U14_Z_5) );
  NOR2_X2 U109 ( .A1(n1065), .A2(n1094), .ZN(U11_Z_5) );
  NOR2_X2 U110 ( .A1(n1067), .A2(n1095), .ZN(U8_Z_5) );
  INV_X4 U111 ( .A(divisor[6]), .ZN(n1228) );
  NOR2_X2 U113 ( .A1(n1182), .A2(n1070), .ZN(U20_Z_6) );
  NOR2_X2 U114 ( .A1(n1063), .A2(n1096), .ZN(U17_Z_6) );
  NOR2_X2 U115 ( .A1(n1064), .A2(n1097), .ZN(U14_Z_6) );
  NOR2_X2 U116 ( .A1(n1065), .A2(n1098), .ZN(U11_Z_6) );
  NOR2_X2 U117 ( .A1(n1067), .A2(n1099), .ZN(U8_Z_6) );
  INV_X4 U118 ( .A(divisor[7]), .ZN(n1227) );
  NOR2_X2 U119 ( .A1(n1182), .A2(n1071), .ZN(U20_Z_7) );
  NOR2_X2 U120 ( .A1(n1063), .A2(n1100), .ZN(U17_Z_7) );
  NOR2_X2 U121 ( .A1(n1064), .A2(n1101), .ZN(U14_Z_7) );
  NOR2_X2 U122 ( .A1(n1065), .A2(n1102), .ZN(U11_Z_7) );
  NOR2_X2 U124 ( .A1(n1067), .A2(n1103), .ZN(U8_Z_7) );
  INV_X4 U125 ( .A(divisor[8]), .ZN(n1226) );
  NOR2_X2 U126 ( .A1(n1182), .A2(n1080), .ZN(U20_Z_8) );
  NOR2_X2 U127 ( .A1(n1063), .A2(n1150), .ZN(U17_Z_8) );
  NOR2_X2 U128 ( .A1(n1064), .A2(n1151), .ZN(U14_Z_8) );
  NOR2_X2 U129 ( .A1(n1065), .A2(n1152), .ZN(U11_Z_8) );
  NOR2_X2 U130 ( .A1(n1067), .A2(n1153), .ZN(U8_Z_8) );
  INV_X4 U131 ( .A(divisor[9]), .ZN(n1225) );
  NOR2_X2 U132 ( .A1(n1182), .A2(n1212), .ZN(U20_Z_9) );
  NOR2_X2 U134 ( .A1(n1063), .A2(n1104), .ZN(U17_Z_9) );
  NOR2_X2 U135 ( .A1(n1064), .A2(n1105), .ZN(U14_Z_9) );
  NOR2_X2 U136 ( .A1(n1065), .A2(n1106), .ZN(U11_Z_9) );
  NOR2_X2 U137 ( .A1(n1067), .A2(n1107), .ZN(U8_Z_9) );
  INV_X4 U138 ( .A(divisor[10]), .ZN(n1224) );
  NOR2_X2 U139 ( .A1(n1182), .A2(n1081), .ZN(U20_Z_10) );
  NOR2_X2 U140 ( .A1(n1063), .A2(n1154), .ZN(U17_Z_10) );
  NOR2_X2 U141 ( .A1(n1064), .A2(n1155), .ZN(U14_Z_10) );
  NOR2_X2 U142 ( .A1(n1065), .A2(n1156), .ZN(U11_Z_10) );
  NOR2_X2 U143 ( .A1(n1067), .A2(n1157), .ZN(U8_Z_10) );
  INV_X4 U144 ( .A(divisor[11]), .ZN(n1223) );
  NOR2_X2 U150 ( .A1(n1182), .A2(n1213), .ZN(U20_Z_11) );
  NOR2_X2 U151 ( .A1(n1063), .A2(n1108), .ZN(U17_Z_11) );
  NOR2_X2 U152 ( .A1(n1064), .A2(n1109), .ZN(U14_Z_11) );
  NOR2_X2 U153 ( .A1(n1065), .A2(n1110), .ZN(U11_Z_11) );
  NOR2_X2 U154 ( .A1(n1067), .A2(n1111), .ZN(U8_Z_11) );
  INV_X4 U159 ( .A(divisor[12]), .ZN(n1222) );
  NOR2_X2 U160 ( .A1(n1182), .A2(n1082), .ZN(U20_Z_12) );
  NOR2_X2 U161 ( .A1(n1063), .A2(n1158), .ZN(U17_Z_12) );
  NOR2_X2 U162 ( .A1(n1064), .A2(n1159), .ZN(U14_Z_12) );
  NOR2_X2 U163 ( .A1(n1065), .A2(n1160), .ZN(U11_Z_12) );
  NOR2_X2 U164 ( .A1(n1067), .A2(n1161), .ZN(U8_Z_12) );
  INV_X4 U165 ( .A(divisor[13]), .ZN(n1221) );
  NOR2_X2 U166 ( .A1(n1182), .A2(n1072), .ZN(U20_Z_13) );
  NOR2_X2 U168 ( .A1(n1063), .A2(n1112), .ZN(U17_Z_13) );
  NOR2_X2 U169 ( .A1(n1064), .A2(n1113), .ZN(U14_Z_13) );
  NOR2_X2 U170 ( .A1(n1065), .A2(n1114), .ZN(U11_Z_13) );
  NOR2_X2 U171 ( .A1(n1067), .A2(n1115), .ZN(U8_Z_13) );
  INV_X4 U172 ( .A(divisor[14]), .ZN(n1220) );
  NOR2_X2 U173 ( .A1(n1182), .A2(n1073), .ZN(U20_Z_14) );
  NOR2_X2 U174 ( .A1(n1063), .A2(n1116), .ZN(U17_Z_14) );
  NOR2_X2 U175 ( .A1(n1064), .A2(n1117), .ZN(U14_Z_14) );
  NOR2_X2 U176 ( .A1(n1065), .A2(n1118), .ZN(U11_Z_14) );
  NOR2_X2 U177 ( .A1(n1067), .A2(n1119), .ZN(U8_Z_14) );
  INV_X4 U179 ( .A(divisor[15]), .ZN(n1219) );
  NOR2_X2 U180 ( .A1(n1182), .A2(n1074), .ZN(U20_Z_15) );
  NOR2_X2 U181 ( .A1(n1063), .A2(n1120), .ZN(U17_Z_15) );
  NOR2_X2 U182 ( .A1(n1064), .A2(n1121), .ZN(U14_Z_15) );
  NOR2_X2 U183 ( .A1(n1065), .A2(n1122), .ZN(U11_Z_15) );
  NOR2_X2 U188 ( .A1(n1067), .A2(n1123), .ZN(U8_Z_15) );
  INV_X4 U189 ( .A(divisor[16]), .ZN(n1218) );
  NOR2_X2 U190 ( .A1(n1182), .A2(n1083), .ZN(U20_Z_16) );
  NOR2_X2 U191 ( .A1(n1063), .A2(n1214), .ZN(U17_Z_16) );
  NOR2_X2 U192 ( .A1(n1064), .A2(n1162), .ZN(U14_Z_16) );
  NOR2_X2 U193 ( .A1(n1065), .A2(n1163), .ZN(U11_Z_16) );
  NOR2_X2 U194 ( .A1(n1067), .A2(n1164), .ZN(U8_Z_16) );
  INV_X4 U195 ( .A(divisor[17]), .ZN(n1217) );
  NOR2_X2 U197 ( .A1(n1182), .A2(n1075), .ZN(U20_Z_17) );
  NOR2_X2 U198 ( .A1(n1063), .A2(n1124), .ZN(U17_Z_17) );
  NOR2_X2 U199 ( .A1(n1064), .A2(n1125), .ZN(U14_Z_17) );
  NOR2_X2 U200 ( .A1(n1065), .A2(n1126), .ZN(U11_Z_17) );
  INV_X4 U201 ( .A(divisor[18]), .ZN(n1216) );
  NOR2_X2 U202 ( .A1(n1182), .A2(n1076), .ZN(U20_Z_18) );
  NOR2_X2 U203 ( .A1(n1063), .A2(n1165), .ZN(U17_Z_18) );
  NOR2_X2 U204 ( .A1(n1064), .A2(n1166), .ZN(U14_Z_18) );
  NOR2_X2 U205 ( .A1(n1065), .A2(n1167), .ZN(U11_Z_18) );
  NOR2_X2 U206 ( .A1(n1067), .A2(n1168), .ZN(U8_Z_18) );
  AND2_X1 U208 ( .A1(U9_DATA1_7), .A2(n355), .ZN(U9_Z_7) );
  AND2_X1 U209 ( .A1(U9_DATA1_8), .A2(n355), .ZN(U9_Z_8) );
  AND2_X1 U210 ( .A1(U9_DATA1_9), .A2(n355), .ZN(U9_Z_9) );
  AND2_X1 U211 ( .A1(U9_DATA1_10), .A2(n355), .ZN(U9_Z_10) );
  AND2_X1 U212 ( .A1(U9_DATA1_11), .A2(n355), .ZN(U9_Z_11) );
  AND2_X1 U213 ( .A1(U9_DATA1_12), .A2(n355), .ZN(U9_Z_12) );
  AND2_X1 U214 ( .A1(U9_DATA1_13), .A2(n355), .ZN(U9_Z_13) );
  AND2_X1 U215 ( .A1(U9_DATA1_14), .A2(n355), .ZN(U9_Z_14) );
  AND2_X1 U216 ( .A1(U9_DATA1_15), .A2(n355), .ZN(U9_Z_15) );
  AND2_X1 U218 ( .A1(U9_DATA1_16), .A2(n355), .ZN(U9_Z_16) );
  AND2_X1 U219 ( .A1(U9_DATA1_17), .A2(n355), .ZN(U9_Z_17) );
  AND2_X1 U220 ( .A1(U9_DATA1_18), .A2(n355), .ZN(U9_Z_18) );
  AND2_X1 U221 ( .A1(U9_DATA1_19), .A2(n355), .ZN(U9_Z_19) );
  AND2_X1 U222 ( .A1(U9_DATA1_20), .A2(n355), .ZN(U9_Z_20) );
  AND2_X1 U223 ( .A1(U9_DATA1_21), .A2(n355), .ZN(U9_Z_21) );
  AND2_X1 U224 ( .A1(U9_DATA1_22), .A2(n355), .ZN(U9_Z_22) );
  AND2_X1 U225 ( .A1(U9_DATA1_23), .A2(n355), .ZN(U9_Z_23) );
  AND2_X1 U226 ( .A1(U9_DATA1_24), .A2(n355), .ZN(U9_Z_24) );
  AND2_X1 U227 ( .A1(U9_DATA1_25), .A2(n355), .ZN(U9_Z_25) );
  AND2_X1 U228 ( .A1(U9_DATA1_26), .A2(n355), .ZN(U9_Z_26) );
  AND2_X1 U229 ( .A1(U9_DATA1_27), .A2(n355), .ZN(U9_Z_27) );
  AND2_X1 U230 ( .A1(U12_DATA1_7), .A2(n491), .ZN(U12_Z_7) );
  AND2_X1 U231 ( .A1(U12_DATA1_8), .A2(n491), .ZN(U12_Z_8) );
  AND2_X1 U232 ( .A1(U12_DATA1_9), .A2(n491), .ZN(U12_Z_9) );
  AND2_X1 U233 ( .A1(U12_DATA1_10), .A2(n491), .ZN(U12_Z_10) );
  AND2_X1 U238 ( .A1(U12_DATA1_11), .A2(n491), .ZN(U12_Z_11) );
  AND2_X1 U239 ( .A1(U12_DATA1_12), .A2(n491), .ZN(U12_Z_12) );
  AND2_X1 U240 ( .A1(U12_DATA1_13), .A2(n491), .ZN(U12_Z_13) );
  AND2_X1 U241 ( .A1(U12_DATA1_14), .A2(n491), .ZN(U12_Z_14) );
  AND2_X1 U242 ( .A1(U12_DATA1_15), .A2(n491), .ZN(U12_Z_15) );
  AND2_X1 U243 ( .A1(U12_DATA1_16), .A2(n491), .ZN(U12_Z_16) );
  AND2_X1 U244 ( .A1(U12_DATA1_17), .A2(n491), .ZN(U12_Z_17) );
  AND2_X1 U245 ( .A1(U12_DATA1_18), .A2(n491), .ZN(U12_Z_18) );
  AND2_X1 U247 ( .A1(U12_DATA1_19), .A2(n491), .ZN(U12_Z_19) );
  AND2_X1 U248 ( .A1(U12_DATA1_20), .A2(n491), .ZN(U12_Z_20) );
  AND2_X1 U249 ( .A1(U12_DATA1_21), .A2(n491), .ZN(U12_Z_21) );
  AND2_X1 U250 ( .A1(U12_DATA1_22), .A2(n491), .ZN(U12_Z_22) );
  AND2_X1 U251 ( .A1(U12_DATA1_23), .A2(n491), .ZN(U12_Z_23) );
  AND2_X1 U252 ( .A1(U12_DATA1_24), .A2(n491), .ZN(U12_Z_24) );
  AND2_X1 U253 ( .A1(U12_DATA1_25), .A2(n491), .ZN(U12_Z_25) );
  AND2_X1 U254 ( .A1(U12_DATA1_26), .A2(n491), .ZN(U12_Z_26) );
  AND2_X1 U255 ( .A1(U12_DATA1_27), .A2(n491), .ZN(U12_Z_27) );
  AND2_X1 U256 ( .A1(U15_DATA1_7), .A2(n625), .ZN(U15_Z_7) );
  AND2_X1 U258 ( .A1(U15_DATA1_8), .A2(n625), .ZN(U15_Z_8) );
  AND2_X1 U259 ( .A1(U15_DATA1_9), .A2(n625), .ZN(U15_Z_9) );
  AND2_X1 U260 ( .A1(U15_DATA1_10), .A2(n625), .ZN(U15_Z_10) );
  AND2_X1 U261 ( .A1(U15_DATA1_11), .A2(n625), .ZN(U15_Z_11) );
  AND2_X1 U262 ( .A1(U15_DATA1_12), .A2(n625), .ZN(U15_Z_12) );
  AND2_X1 U263 ( .A1(U15_DATA1_13), .A2(n625), .ZN(U15_Z_13) );
  AND2_X1 U264 ( .A1(U15_DATA1_14), .A2(n625), .ZN(U15_Z_14) );
  AND2_X1 U265 ( .A1(U15_DATA1_15), .A2(n625), .ZN(U15_Z_15) );
  AND2_X1 U266 ( .A1(U15_DATA1_16), .A2(n625), .ZN(U15_Z_16) );
  AND2_X1 U268 ( .A1(U15_DATA1_17), .A2(n625), .ZN(U15_Z_17) );
  AND2_X1 U269 ( .A1(U15_DATA1_18), .A2(n625), .ZN(U15_Z_18) );
  AND2_X1 U270 ( .A1(U15_DATA1_19), .A2(n625), .ZN(U15_Z_19) );
  AND2_X1 U271 ( .A1(U15_DATA1_20), .A2(n625), .ZN(U15_Z_20) );
  AND2_X1 U272 ( .A1(U15_DATA1_21), .A2(n625), .ZN(U15_Z_21) );
  AND2_X1 U273 ( .A1(U15_DATA1_22), .A2(n625), .ZN(U15_Z_22) );
  AND2_X1 U274 ( .A1(U15_DATA1_23), .A2(n625), .ZN(U15_Z_23) );
  AND2_X1 U275 ( .A1(U15_DATA1_24), .A2(n625), .ZN(U15_Z_24) );
  AND2_X1 U276 ( .A1(U15_DATA1_25), .A2(n625), .ZN(U15_Z_25) );
  AND2_X1 U277 ( .A1(U15_DATA1_26), .A2(n625), .ZN(U15_Z_26) );
  AND2_X1 U278 ( .A1(U15_DATA1_27), .A2(n625), .ZN(U15_Z_27) );
  AND2_X1 U280 ( .A1(U18_DATA1_7), .A2(n1068), .ZN(U18_Z_7) );
  AND2_X1 U281 ( .A1(U18_DATA1_8), .A2(n1068), .ZN(U18_Z_8) );
  AND2_X1 U282 ( .A1(U18_DATA1_9), .A2(n1068), .ZN(U18_Z_9) );
  AND2_X1 U283 ( .A1(U18_DATA1_10), .A2(n1068), .ZN(U18_Z_10) );
  AND2_X1 U284 ( .A1(U18_DATA1_11), .A2(n1068), .ZN(U18_Z_11) );
  AND2_X1 U289 ( .A1(U18_DATA1_12), .A2(n1068), .ZN(U18_Z_12) );
  AND2_X1 U290 ( .A1(U18_DATA1_13), .A2(n1068), .ZN(U18_Z_13) );
  AND2_X1 U291 ( .A1(U18_DATA1_14), .A2(n1068), .ZN(U18_Z_14) );
  AND2_X1 U292 ( .A1(U18_DATA1_15), .A2(n1068), .ZN(U18_Z_15) );
  AND2_X1 U293 ( .A1(U18_DATA1_16), .A2(n1068), .ZN(U18_Z_16) );
  AND2_X1 U294 ( .A1(U18_DATA1_17), .A2(n1068), .ZN(U18_Z_17) );
  AND2_X1 U295 ( .A1(U18_DATA1_18), .A2(n1068), .ZN(U18_Z_18) );
  AND2_X1 U296 ( .A1(U18_DATA1_19), .A2(n1068), .ZN(U18_Z_19) );
  AND2_X1 U298 ( .A1(U18_DATA1_20), .A2(n1068), .ZN(U18_Z_20) );
  AND2_X1 U299 ( .A1(U18_DATA1_21), .A2(n1068), .ZN(U18_Z_21) );
  AND2_X1 U300 ( .A1(U18_DATA1_22), .A2(n1068), .ZN(U18_Z_22) );
  AND2_X1 U301 ( .A1(U18_DATA1_23), .A2(n1068), .ZN(U18_Z_23) );
  AND2_X1 U302 ( .A1(U18_DATA1_24), .A2(n1068), .ZN(U18_Z_24) );
  AND2_X1 U303 ( .A1(U18_DATA1_25), .A2(n1068), .ZN(U18_Z_25) );
  AND2_X1 U304 ( .A1(U18_DATA1_26), .A2(n1068), .ZN(U18_Z_26) );
  AND2_X1 U305 ( .A1(U18_DATA1_27), .A2(n1068), .ZN(U18_Z_27) );
  AND2_X1 U306 ( .A1(U21_DATA1_7), .A2(n887), .ZN(U21_Z_7) );
  AND2_X1 U307 ( .A1(U21_DATA1_8), .A2(n887), .ZN(U21_Z_8) );
  AND2_X1 U309 ( .A1(U21_DATA1_9), .A2(n887), .ZN(U21_Z_9) );
  AND2_X1 U310 ( .A1(U21_DATA1_10), .A2(n887), .ZN(U21_Z_10) );
  AND2_X1 U311 ( .A1(U21_DATA1_11), .A2(n887), .ZN(U21_Z_11) );
  AND2_X1 U312 ( .A1(U21_DATA1_12), .A2(n887), .ZN(U21_Z_12) );
  AND2_X1 U313 ( .A1(U21_DATA1_13), .A2(n887), .ZN(U21_Z_13) );
  AND2_X1 U314 ( .A1(U21_DATA1_14), .A2(n887), .ZN(U21_Z_14) );
  AND2_X1 U315 ( .A1(U21_DATA1_15), .A2(n887), .ZN(U21_Z_15) );
  AND2_X1 U316 ( .A1(U21_DATA1_16), .A2(n887), .ZN(U21_Z_16) );
  AND2_X1 U317 ( .A1(U21_DATA1_17), .A2(n887), .ZN(U21_Z_17) );
  AND2_X1 U319 ( .A1(U21_DATA1_18), .A2(n887), .ZN(U21_Z_18) );
  AND2_X1 U320 ( .A1(U21_DATA1_19), .A2(n887), .ZN(U21_Z_19) );
  AND2_X1 U321 ( .A1(U21_DATA1_20), .A2(n887), .ZN(U21_Z_20) );
  AND2_X1 U322 ( .A1(U21_DATA1_21), .A2(n887), .ZN(U21_Z_21) );
  AND2_X1 U323 ( .A1(U21_DATA1_22), .A2(n887), .ZN(U21_Z_22) );
  AND2_X1 U324 ( .A1(U21_DATA1_23), .A2(n887), .ZN(U21_Z_23) );
  AND2_X1 U325 ( .A1(U21_DATA1_24), .A2(n887), .ZN(U21_Z_24) );
  AND2_X1 U326 ( .A1(U21_DATA1_25), .A2(n887), .ZN(U21_Z_25) );
  AND2_X1 U327 ( .A1(U21_DATA1_26), .A2(n887), .ZN(U21_Z_26) );
  AND2_X1 U328 ( .A1(U21_DATA1_27), .A2(n887), .ZN(U21_Z_27) );
  AND2_X1 U329 ( .A1(U24_DATA1_7), .A2(n1183), .ZN(U24_Z_7) );
  AND2_X1 U332 ( .A1(U24_DATA1_8), .A2(start), .ZN(U24_Z_8) );
  AND2_X1 U333 ( .A1(U24_DATA1_9), .A2(n1183), .ZN(U24_Z_9) );
  AND2_X1 U334 ( .A1(U24_DATA1_10), .A2(start), .ZN(U24_Z_10) );
  AND2_X1 U335 ( .A1(U24_DATA1_11), .A2(n1183), .ZN(U24_Z_11) );
  AND2_X1 U336 ( .A1(U24_DATA1_12), .A2(start), .ZN(U24_Z_12) );
  AND2_X1 U341 ( .A1(U24_DATA1_13), .A2(n1183), .ZN(U24_Z_13) );
  AND2_X1 U342 ( .A1(U24_DATA1_14), .A2(start), .ZN(U24_Z_14) );
  AND2_X1 U343 ( .A1(U24_DATA1_15), .A2(start), .ZN(U24_Z_15) );
  AND2_X1 U344 ( .A1(U24_DATA1_16), .A2(start), .ZN(U24_Z_16) );
  AND2_X1 U345 ( .A1(U24_DATA1_17), .A2(start), .ZN(U24_Z_17) );
  AND2_X1 U346 ( .A1(U24_DATA1_18), .A2(start), .ZN(U24_Z_18) );
  AND2_X1 U347 ( .A1(U24_DATA1_19), .A2(start), .ZN(U24_Z_19) );
  AND2_X1 U348 ( .A1(U24_DATA1_20), .A2(start), .ZN(U24_Z_20) );
  AND2_X1 U350 ( .A1(U24_DATA1_21), .A2(start), .ZN(U24_Z_21) );
  AND2_X1 U351 ( .A1(U24_DATA1_22), .A2(n1183), .ZN(U24_Z_22) );
  AND2_X1 U352 ( .A1(U24_DATA1_23), .A2(n1183), .ZN(U24_Z_23) );
  AND2_X1 U353 ( .A1(U24_DATA1_24), .A2(n1183), .ZN(U24_Z_24) );
  AND2_X1 U354 ( .A1(U24_DATA1_25), .A2(n1183), .ZN(U24_Z_25) );
  AND2_X1 U355 ( .A1(U24_DATA1_26), .A2(n1183), .ZN(U24_Z_26) );
  AND2_X1 U356 ( .A1(U24_DATA1_27), .A2(n1183), .ZN(U24_Z_27) );
  AND2_X1 U357 ( .A1(U6_DATA1_27), .A2(n217), .ZN(U6_Z_27) );
  AND2_X1 U358 ( .A1(U6_DATA1_26), .A2(n217), .ZN(U6_Z_26) );
  AND2_X1 U359 ( .A1(U6_DATA1_25), .A2(n217), .ZN(U6_Z_25) );
  AND2_X1 U361 ( .A1(U6_DATA1_24), .A2(n217), .ZN(U6_Z_24) );
  AND2_X1 U362 ( .A1(U6_DATA1_23), .A2(n217), .ZN(U6_Z_23) );
  AND2_X1 U363 ( .A1(U6_DATA1_22), .A2(n217), .ZN(U6_Z_22) );
  AND2_X1 U364 ( .A1(U6_DATA1_21), .A2(n217), .ZN(U6_Z_21) );
  AND2_X1 U365 ( .A1(U6_DATA1_20), .A2(n217), .ZN(U6_Z_20) );
  AND2_X1 U366 ( .A1(U6_DATA1_19), .A2(n217), .ZN(U6_Z_19) );
  AND2_X1 U367 ( .A1(U6_DATA1_18), .A2(n217), .ZN(U6_Z_18) );
  AND2_X1 U368 ( .A1(U6_DATA1_17), .A2(n217), .ZN(U6_Z_17) );
  AND2_X1 U369 ( .A1(U6_DATA1_16), .A2(n217), .ZN(U6_Z_16) );
  AND2_X1 U371 ( .A1(U6_DATA1_15), .A2(n217), .ZN(U6_Z_15) );
  AND2_X1 U372 ( .A1(U6_DATA1_14), .A2(n217), .ZN(U6_Z_14) );
  AND2_X1 U373 ( .A1(U6_DATA1_13), .A2(n217), .ZN(U6_Z_13) );
  AND2_X1 U374 ( .A1(U6_DATA1_12), .A2(n217), .ZN(U6_Z_12) );
  AND2_X1 U375 ( .A1(U6_DATA1_11), .A2(n217), .ZN(U6_Z_11) );
  AND2_X1 U376 ( .A1(U6_DATA1_10), .A2(n217), .ZN(U6_Z_10) );
  AND2_X1 U377 ( .A1(U6_DATA1_9), .A2(n217), .ZN(U6_Z_9) );
  AND2_X1 U378 ( .A1(U6_DATA1_8), .A2(n217), .ZN(U6_Z_8) );
  NOR2_X2 U379 ( .A1(n1066), .A2(n1169), .ZN(U5_Z_18) );
  NOR2_X2 U380 ( .A1(n1066), .A2(n1215), .ZN(U5_Z_17) );
  NOR2_X2 U381 ( .A1(n1066), .A2(n1170), .ZN(U5_Z_16) );
  NOR2_X2 U385 ( .A1(n1066), .A2(n1127), .ZN(U5_Z_15) );
  NOR2_X2 U386 ( .A1(n1066), .A2(n1128), .ZN(U5_Z_14) );
  NOR2_X2 U387 ( .A1(n1066), .A2(n1129), .ZN(U5_Z_13) );
  NOR2_X2 U388 ( .A1(n1066), .A2(n1171), .ZN(U5_Z_12) );
  NOR2_X2 U389 ( .A1(n1066), .A2(n1130), .ZN(U5_Z_11) );
  NOR2_X2 U390 ( .A1(n1066), .A2(n1172), .ZN(U5_Z_10) );
  NOR2_X2 U391 ( .A1(n1066), .A2(n1131), .ZN(U5_Z_9) );
  NOR2_X2 U392 ( .A1(n1066), .A2(n1173), .ZN(U5_Z_8) );
  NOR2_X2 U393 ( .A1(n1066), .A2(n1132), .ZN(U5_Z_7) );
  NOR2_X2 U394 ( .A1(n1066), .A2(n1133), .ZN(U5_Z_6) );
  NOR2_X2 U395 ( .A1(n1066), .A2(n1134), .ZN(U5_Z_5) );
  NOR2_X2 U396 ( .A1(n1066), .A2(n1174), .ZN(U5_Z_4) );
  NOR2_X2 U397 ( .A1(n1066), .A2(n1135), .ZN(U5_Z_3) );
  NOR2_X2 U398 ( .A1(n1066), .A2(n1175), .ZN(U5_Z_2) );
  NOR2_X2 U399 ( .A1(n1066), .A2(n1136), .ZN(U5_Z_1) );
  NOR2_X2 U400 ( .A1(n1066), .A2(n1141), .ZN(U5_Z_0) );
  AND2_X1 U401 ( .A1(U4_DATA1_0), .A2(n217), .ZN(U4_Z_0) );
  AND2_X1 U402 ( .A1(U7_DATA1_0), .A2(n355), .ZN(U7_Z_0) );
  AND2_X1 U403 ( .A1(U4_DATA1_1), .A2(n217), .ZN(U4_Z_1) );
  AND2_X1 U404 ( .A1(U10_DATA1_0), .A2(n491), .ZN(U10_Z_0) );
  AND2_X1 U405 ( .A1(U7_DATA1_1), .A2(n355), .ZN(U7_Z_1) );
  AND2_X1 U406 ( .A1(U13_DATA1_0), .A2(n625), .ZN(U13_Z_0) );
  AND2_X1 U407 ( .A1(U10_DATA1_1), .A2(n491), .ZN(U10_Z_1) );
  AND2_X1 U408 ( .A1(U16_DATA1_0), .A2(n1068), .ZN(U16_Z_0) );
  AND2_X1 U409 ( .A1(U13_DATA1_1), .A2(n625), .ZN(U13_Z_1) );
  AND2_X1 U410 ( .A1(U19_DATA1_0), .A2(n887), .ZN(U19_Z_0) );
  AND2_X1 U411 ( .A1(U16_DATA1_1), .A2(n1068), .ZN(U16_Z_1) );
  AND2_X1 U412 ( .A1(U22_DATA1_0), .A2(n1183), .ZN(U22_Z_0) );
  AND2_X1 U413 ( .A1(U19_DATA1_1), .A2(n887), .ZN(U19_Z_1) );
  BUF_X8 U28 ( .A(reset_n), .Z(n1189) );
endmodule


module Output_Result ( clock, reset_n, DataIn, StartIn, Divisor, StartOut, 
        DataOut );
  input [27:0] DataIn;
  input [19:0] Divisor;
  output [7:0] DataOut;
  input clock, reset_n, StartIn;
  output StartOut;


  pipeline_divider divider ( .clock(clock), .reset_n(reset_n), .start(StartIn), 
        .divided(DataIn), .divisor(Divisor), .q(DataOut), .StartOut(StartOut)
         );
endmodule


module Output_Store ( clock, reset_n, StartIn, ResultIn, WriteBus, 
        WriteAddress, WriteEnable, output_base_offset );
  input [7:0] ResultIn;
  output [127:0] WriteBus;
  output [15:0] WriteAddress;
  input clock, reset_n, StartIn, output_base_offset;
  output WriteEnable;
  wire   U5_DATA1_0, U5_DATA1_1, U5_DATA1_2, U5_DATA1_3, U5_DATA1_4,
         U5_DATA1_5, U5_DATA1_6, U5_DATA1_7, U5_DATA1_8, U5_DATA1_9,
         U5_DATA1_10, U5_DATA1_11, U5_DATA1_12, U5_DATA1_13, U5_DATA1_14,
         U5_DATA1_15, U5_DATA1_16, U5_DATA1_17, U5_DATA1_18, U5_DATA1_19,
         U5_DATA1_20, U5_DATA1_21, U5_DATA1_22, U5_DATA1_23, U5_DATA1_24,
         U5_DATA1_25, U5_DATA1_26, U5_DATA1_27, U5_DATA1_28, U5_DATA1_29,
         U5_DATA1_30, U5_DATA1_31, U5_DATA1_32, U5_DATA1_33, U5_DATA1_34,
         U5_DATA1_35, U5_DATA1_36, U5_DATA1_37, U5_DATA1_38, U5_DATA1_39,
         U5_DATA1_40, U5_DATA1_41, U5_DATA1_42, U5_DATA1_43, U5_DATA1_44,
         U5_DATA1_45, U5_DATA1_46, U5_DATA1_47, U5_DATA1_48, U5_DATA1_49,
         U5_DATA1_50, U5_DATA1_51, U5_DATA1_52, U5_DATA1_53, U5_DATA1_54,
         U5_DATA1_55, U5_DATA1_56, U5_DATA1_57, U5_DATA1_58, U5_DATA1_59,
         U5_DATA1_60, U5_DATA1_61, U5_DATA1_62, U5_DATA1_63, U5_DATA1_64,
         U5_DATA1_65, U5_DATA1_66, U5_DATA1_67, U5_DATA1_68, U5_DATA1_69,
         U5_DATA1_70, U5_DATA1_71, U5_DATA1_72, U5_DATA1_73, U5_DATA1_74,
         U5_DATA1_75, U5_DATA1_76, U5_DATA1_77, U5_DATA1_78, U5_DATA1_79,
         U5_DATA1_80, U5_DATA1_81, U5_DATA1_82, U5_DATA1_83, U5_DATA1_84,
         U5_DATA1_85, U5_DATA1_86, U5_DATA1_87, U5_DATA1_88, U5_DATA1_89,
         U5_DATA1_90, U5_DATA1_91, U5_DATA1_92, U5_DATA1_93, U5_DATA1_94,
         U5_DATA1_95, U5_DATA1_96, U5_DATA1_97, U5_DATA1_98, U5_DATA1_99,
         U5_DATA1_100, U5_DATA1_101, U5_DATA1_102, U5_DATA1_103, U5_DATA1_104,
         U5_DATA1_105, U5_DATA1_106, U5_DATA1_107, U5_DATA1_108, U5_DATA1_109,
         U5_DATA1_110, U5_DATA1_111, U5_DATA1_112, U5_DATA1_113, U5_DATA1_114,
         U5_DATA1_115, U5_DATA1_116, U5_DATA1_117, U5_DATA1_118, U5_DATA1_119,
         U5_DATA1_120, U5_DATA1_121, U5_DATA1_122, U5_DATA1_123, U5_DATA1_124,
         U5_DATA1_125, U5_DATA1_126, U5_DATA1_127, U4_Z_0, U4_Z_1, U4_Z_2,
         U4_Z_3, U4_DATA2_1, U4_DATA2_2, U4_DATA2_3, U4_DATA2_4,
         sub_46_carry_2_, sub_46_carry_3_, sub_46_A_0_, sub_46_A_1_,
         sub_46_A_2_, sub_46_A_3_, sub_46_A_4_, add_37_A_0_, add_37_A_1_,
         add_37_A_2_, add_37_A_3_, add_37_A_4_, add_37_A_5_, add_37_A_6_,
         add_37_A_7_, add_37_A_8_, add_37_A_9_, add_37_A_10_, add_37_A_11_,
         add_37_A_12_, add_37_A_13_, add_37_A_14_, add_37_A_15_, n146, n147,
         n148, n149, n151, n155, n177, n180, n181, n182, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823;

  XNOR2_X2 sub_46_U1_A_1 ( .A(sub_46_A_1_), .B(sub_46_A_0_), .ZN(U4_DATA2_1)
         );
  OR2_X1 sub_46_U1_B_1 ( .A1(sub_46_A_1_), .A2(sub_46_A_0_), .ZN(
        sub_46_carry_2_) );
  XNOR2_X2 sub_46_U1_A_2 ( .A(sub_46_A_2_), .B(sub_46_carry_2_), .ZN(
        U4_DATA2_2) );
  OR2_X1 sub_46_U1_B_2 ( .A1(sub_46_A_2_), .A2(sub_46_carry_2_), .ZN(
        sub_46_carry_3_) );
  XNOR2_X2 sub_46_U1_A_3 ( .A(sub_46_A_3_), .B(sub_46_carry_3_), .ZN(
        U4_DATA2_3) );
  DFFS_X2 short_count_reg_0_ ( .D(U4_Z_0), .CK(clock), .SN(n738), .Q(
        sub_46_A_0_), .QN(n148) );
  DFFS_X2 short_count_reg_1_ ( .D(U4_Z_1), .CK(clock), .SN(n737), .Q(
        sub_46_A_1_) );
  DFFS_X2 short_count_reg_2_ ( .D(U4_Z_2), .CK(clock), .SN(n737), .Q(
        sub_46_A_2_), .QN(n147) );
  DFFS_X2 short_count_reg_3_ ( .D(U4_Z_3), .CK(clock), .SN(n738), .Q(
        sub_46_A_3_), .QN(n146) );
  SDFFR_X2 short_count_reg_4_ ( .D(1'b0), .SI(n808), .SE(U4_DATA2_4), .CK(
        clock), .RN(n738), .Q(sub_46_A_4_) );
  NOR2_X2 U161 ( .A1(n146), .A2(sub_46_A_4_), .ZN(n177) );
  NAND2_X2 U172 ( .A1(sub_46_A_0_), .A2(n808), .ZN(U4_Z_0) );
  NOR2_X2 U177 ( .A1(sub_46_A_3_), .A2(sub_46_A_4_), .ZN(n180) );
  OR2_X1 U196 ( .A1(U4_DATA2_3), .A2(n155), .ZN(U4_Z_3) );
  OR2_X1 U197 ( .A1(U4_DATA2_2), .A2(n155), .ZN(U4_Z_2) );
  OR2_X1 U198 ( .A1(U4_DATA2_1), .A2(n155), .ZN(U4_Z_1) );
  DLH_X2 data_reg_127_ ( .G(n584), .D(ResultIn[7]), .Q(U5_DATA1_127) );
  DLH_X2 data_reg_126_ ( .G(n584), .D(ResultIn[6]), .Q(U5_DATA1_126) );
  DLH_X2 data_reg_125_ ( .G(n584), .D(ResultIn[5]), .Q(U5_DATA1_125) );
  DLH_X2 data_reg_124_ ( .G(n584), .D(ResultIn[4]), .Q(U5_DATA1_124) );
  DLH_X2 data_reg_123_ ( .G(n584), .D(ResultIn[3]), .Q(U5_DATA1_123) );
  DLH_X2 data_reg_122_ ( .G(n584), .D(ResultIn[2]), .Q(U5_DATA1_122) );
  DLH_X2 data_reg_121_ ( .G(n584), .D(ResultIn[1]), .Q(U5_DATA1_121) );
  DLH_X2 data_reg_120_ ( .G(n584), .D(ResultIn[0]), .Q(U5_DATA1_120) );
  DLH_X2 data_reg_119_ ( .G(n583), .D(ResultIn[7]), .Q(U5_DATA1_119) );
  DLH_X2 data_reg_118_ ( .G(n583), .D(ResultIn[6]), .Q(U5_DATA1_118) );
  DLH_X2 data_reg_117_ ( .G(n583), .D(ResultIn[5]), .Q(U5_DATA1_117) );
  DLH_X2 data_reg_116_ ( .G(n583), .D(ResultIn[4]), .Q(U5_DATA1_116) );
  DLH_X2 data_reg_115_ ( .G(n583), .D(ResultIn[3]), .Q(U5_DATA1_115) );
  DLH_X2 data_reg_114_ ( .G(n583), .D(ResultIn[2]), .Q(U5_DATA1_114) );
  DLH_X2 data_reg_113_ ( .G(n583), .D(ResultIn[1]), .Q(U5_DATA1_113) );
  DLH_X2 data_reg_112_ ( .G(n583), .D(ResultIn[0]), .Q(U5_DATA1_112) );
  DLH_X2 data_reg_111_ ( .G(n582), .D(ResultIn[7]), .Q(U5_DATA1_111) );
  DLH_X2 data_reg_110_ ( .G(n582), .D(ResultIn[6]), .Q(U5_DATA1_110) );
  DLH_X2 data_reg_109_ ( .G(n582), .D(ResultIn[5]), .Q(U5_DATA1_109) );
  DLH_X2 data_reg_108_ ( .G(n582), .D(ResultIn[4]), .Q(U5_DATA1_108) );
  DLH_X2 data_reg_107_ ( .G(n582), .D(ResultIn[3]), .Q(U5_DATA1_107) );
  DLH_X2 data_reg_106_ ( .G(n582), .D(ResultIn[2]), .Q(U5_DATA1_106) );
  DLH_X2 data_reg_105_ ( .G(n582), .D(ResultIn[1]), .Q(U5_DATA1_105) );
  DLH_X2 data_reg_104_ ( .G(n582), .D(ResultIn[0]), .Q(U5_DATA1_104) );
  DLH_X2 data_reg_103_ ( .G(n581), .D(ResultIn[7]), .Q(U5_DATA1_103) );
  DLH_X2 data_reg_102_ ( .G(n581), .D(ResultIn[6]), .Q(U5_DATA1_102) );
  DLH_X2 data_reg_101_ ( .G(n581), .D(ResultIn[5]), .Q(U5_DATA1_101) );
  DLH_X2 data_reg_100_ ( .G(n581), .D(ResultIn[4]), .Q(U5_DATA1_100) );
  DLH_X2 data_reg_99_ ( .G(n581), .D(ResultIn[3]), .Q(U5_DATA1_99) );
  DLH_X2 data_reg_98_ ( .G(n581), .D(ResultIn[2]), .Q(U5_DATA1_98) );
  DLH_X2 data_reg_97_ ( .G(n581), .D(ResultIn[1]), .Q(U5_DATA1_97) );
  DLH_X2 data_reg_96_ ( .G(n581), .D(ResultIn[0]), .Q(U5_DATA1_96) );
  DLH_X2 data_reg_95_ ( .G(n580), .D(ResultIn[7]), .Q(U5_DATA1_95) );
  DLH_X2 data_reg_94_ ( .G(n580), .D(ResultIn[6]), .Q(U5_DATA1_94) );
  DLH_X2 data_reg_93_ ( .G(n580), .D(ResultIn[5]), .Q(U5_DATA1_93) );
  DLH_X2 data_reg_92_ ( .G(n580), .D(ResultIn[4]), .Q(U5_DATA1_92) );
  DLH_X2 data_reg_91_ ( .G(n580), .D(ResultIn[3]), .Q(U5_DATA1_91) );
  DLH_X2 data_reg_90_ ( .G(n580), .D(ResultIn[2]), .Q(U5_DATA1_90) );
  DLH_X2 data_reg_89_ ( .G(n580), .D(ResultIn[1]), .Q(U5_DATA1_89) );
  DLH_X2 data_reg_88_ ( .G(n580), .D(ResultIn[0]), .Q(U5_DATA1_88) );
  DLH_X2 data_reg_87_ ( .G(n579), .D(ResultIn[7]), .Q(U5_DATA1_87) );
  DLH_X2 data_reg_86_ ( .G(n579), .D(ResultIn[6]), .Q(U5_DATA1_86) );
  DLH_X2 data_reg_85_ ( .G(n579), .D(ResultIn[5]), .Q(U5_DATA1_85) );
  DLH_X2 data_reg_84_ ( .G(n579), .D(ResultIn[4]), .Q(U5_DATA1_84) );
  DLH_X2 data_reg_83_ ( .G(n579), .D(ResultIn[3]), .Q(U5_DATA1_83) );
  DLH_X2 data_reg_82_ ( .G(n579), .D(ResultIn[2]), .Q(U5_DATA1_82) );
  DLH_X2 data_reg_81_ ( .G(n579), .D(ResultIn[1]), .Q(U5_DATA1_81) );
  DLH_X2 data_reg_80_ ( .G(n579), .D(ResultIn[0]), .Q(U5_DATA1_80) );
  DLH_X2 data_reg_79_ ( .G(n725), .D(ResultIn[7]), .Q(U5_DATA1_79) );
  DLH_X2 data_reg_78_ ( .G(n725), .D(ResultIn[6]), .Q(U5_DATA1_78) );
  DLH_X2 data_reg_77_ ( .G(n725), .D(ResultIn[5]), .Q(U5_DATA1_77) );
  DLH_X2 data_reg_76_ ( .G(n725), .D(ResultIn[4]), .Q(U5_DATA1_76) );
  DLH_X2 data_reg_75_ ( .G(n725), .D(ResultIn[3]), .Q(U5_DATA1_75) );
  DLH_X2 data_reg_74_ ( .G(n725), .D(ResultIn[2]), .Q(U5_DATA1_74) );
  DLH_X2 data_reg_73_ ( .G(n725), .D(ResultIn[1]), .Q(U5_DATA1_73) );
  DLH_X2 data_reg_72_ ( .G(n725), .D(ResultIn[0]), .Q(U5_DATA1_72) );
  DLH_X2 data_reg_71_ ( .G(n724), .D(ResultIn[7]), .Q(U5_DATA1_71) );
  DLH_X2 data_reg_70_ ( .G(n724), .D(ResultIn[6]), .Q(U5_DATA1_70) );
  DLH_X2 data_reg_69_ ( .G(n724), .D(ResultIn[5]), .Q(U5_DATA1_69) );
  DLH_X2 data_reg_68_ ( .G(n724), .D(ResultIn[4]), .Q(U5_DATA1_68) );
  DLH_X2 data_reg_67_ ( .G(n724), .D(ResultIn[3]), .Q(U5_DATA1_67) );
  DLH_X2 data_reg_66_ ( .G(n724), .D(ResultIn[2]), .Q(U5_DATA1_66) );
  DLH_X2 data_reg_65_ ( .G(n724), .D(ResultIn[1]), .Q(U5_DATA1_65) );
  DLH_X2 data_reg_64_ ( .G(n724), .D(ResultIn[0]), .Q(U5_DATA1_64) );
  DLH_X2 data_reg_63_ ( .G(n589), .D(ResultIn[7]), .Q(U5_DATA1_63) );
  DLH_X2 data_reg_62_ ( .G(n589), .D(ResultIn[6]), .Q(U5_DATA1_62) );
  DLH_X2 data_reg_61_ ( .G(n589), .D(ResultIn[5]), .Q(U5_DATA1_61) );
  DLH_X2 data_reg_60_ ( .G(n589), .D(ResultIn[4]), .Q(U5_DATA1_60) );
  DLH_X2 data_reg_59_ ( .G(n589), .D(ResultIn[3]), .Q(U5_DATA1_59) );
  DLH_X2 data_reg_58_ ( .G(n589), .D(ResultIn[2]), .Q(U5_DATA1_58) );
  DLH_X2 data_reg_57_ ( .G(n589), .D(ResultIn[1]), .Q(U5_DATA1_57) );
  DLH_X2 data_reg_56_ ( .G(n589), .D(ResultIn[0]), .Q(U5_DATA1_56) );
  DLH_X2 data_reg_55_ ( .G(n723), .D(ResultIn[7]), .Q(U5_DATA1_55) );
  DLH_X2 data_reg_54_ ( .G(n723), .D(ResultIn[6]), .Q(U5_DATA1_54) );
  DLH_X2 data_reg_53_ ( .G(n723), .D(ResultIn[5]), .Q(U5_DATA1_53) );
  DLH_X2 data_reg_52_ ( .G(n723), .D(ResultIn[4]), .Q(U5_DATA1_52) );
  DLH_X2 data_reg_51_ ( .G(n723), .D(ResultIn[3]), .Q(U5_DATA1_51) );
  DLH_X2 data_reg_50_ ( .G(n723), .D(ResultIn[2]), .Q(U5_DATA1_50) );
  DLH_X2 data_reg_49_ ( .G(n723), .D(ResultIn[1]), .Q(U5_DATA1_49) );
  DLH_X2 data_reg_48_ ( .G(n723), .D(ResultIn[0]), .Q(U5_DATA1_48) );
  DLH_X2 data_reg_47_ ( .G(n588), .D(ResultIn[7]), .Q(U5_DATA1_47) );
  DLH_X2 data_reg_46_ ( .G(n588), .D(ResultIn[6]), .Q(U5_DATA1_46) );
  DLH_X2 data_reg_45_ ( .G(n588), .D(ResultIn[5]), .Q(U5_DATA1_45) );
  DLH_X2 data_reg_44_ ( .G(n588), .D(ResultIn[4]), .Q(U5_DATA1_44) );
  DLH_X2 data_reg_43_ ( .G(n588), .D(ResultIn[3]), .Q(U5_DATA1_43) );
  DLH_X2 data_reg_42_ ( .G(n588), .D(ResultIn[2]), .Q(U5_DATA1_42) );
  DLH_X2 data_reg_41_ ( .G(n588), .D(ResultIn[1]), .Q(U5_DATA1_41) );
  DLH_X2 data_reg_40_ ( .G(n588), .D(ResultIn[0]), .Q(U5_DATA1_40) );
  DLH_X2 data_reg_39_ ( .G(n722), .D(ResultIn[7]), .Q(U5_DATA1_39) );
  DLH_X2 data_reg_38_ ( .G(n722), .D(ResultIn[6]), .Q(U5_DATA1_38) );
  DLH_X2 data_reg_37_ ( .G(n722), .D(ResultIn[5]), .Q(U5_DATA1_37) );
  DLH_X2 data_reg_36_ ( .G(n722), .D(ResultIn[4]), .Q(U5_DATA1_36) );
  DLH_X2 data_reg_35_ ( .G(n722), .D(ResultIn[3]), .Q(U5_DATA1_35) );
  DLH_X2 data_reg_34_ ( .G(n722), .D(ResultIn[2]), .Q(U5_DATA1_34) );
  DLH_X2 data_reg_33_ ( .G(n722), .D(ResultIn[1]), .Q(U5_DATA1_33) );
  DLH_X2 data_reg_32_ ( .G(n722), .D(ResultIn[0]), .Q(U5_DATA1_32) );
  DLH_X2 data_reg_31_ ( .G(n587), .D(ResultIn[7]), .Q(U5_DATA1_31) );
  DLH_X2 data_reg_30_ ( .G(n587), .D(ResultIn[6]), .Q(U5_DATA1_30) );
  DLH_X2 data_reg_29_ ( .G(n587), .D(ResultIn[5]), .Q(U5_DATA1_29) );
  DLH_X2 data_reg_28_ ( .G(n587), .D(ResultIn[4]), .Q(U5_DATA1_28) );
  DLH_X2 data_reg_27_ ( .G(n587), .D(ResultIn[3]), .Q(U5_DATA1_27) );
  DLH_X2 data_reg_26_ ( .G(n587), .D(ResultIn[2]), .Q(U5_DATA1_26) );
  DLH_X2 data_reg_25_ ( .G(n587), .D(ResultIn[1]), .Q(U5_DATA1_25) );
  DLH_X2 data_reg_24_ ( .G(n587), .D(ResultIn[0]), .Q(U5_DATA1_24) );
  DLH_X2 data_reg_23_ ( .G(n721), .D(ResultIn[7]), .Q(U5_DATA1_23) );
  DLH_X2 data_reg_22_ ( .G(n721), .D(ResultIn[6]), .Q(U5_DATA1_22) );
  DLH_X2 data_reg_21_ ( .G(n721), .D(ResultIn[5]), .Q(U5_DATA1_21) );
  DLH_X2 data_reg_20_ ( .G(n721), .D(ResultIn[4]), .Q(U5_DATA1_20) );
  DLH_X2 data_reg_19_ ( .G(n721), .D(ResultIn[3]), .Q(U5_DATA1_19) );
  DLH_X2 data_reg_18_ ( .G(n721), .D(ResultIn[2]), .Q(U5_DATA1_18) );
  DLH_X2 data_reg_17_ ( .G(n721), .D(ResultIn[1]), .Q(U5_DATA1_17) );
  DLH_X2 data_reg_16_ ( .G(n721), .D(ResultIn[0]), .Q(U5_DATA1_16) );
  DLH_X2 data_reg_15_ ( .G(n720), .D(ResultIn[7]), .Q(U5_DATA1_15) );
  DLH_X2 data_reg_14_ ( .G(n720), .D(ResultIn[6]), .Q(U5_DATA1_14) );
  DLH_X2 data_reg_13_ ( .G(n720), .D(ResultIn[5]), .Q(U5_DATA1_13) );
  DLH_X2 data_reg_12_ ( .G(n720), .D(ResultIn[4]), .Q(U5_DATA1_12) );
  DLH_X2 data_reg_11_ ( .G(n720), .D(ResultIn[3]), .Q(U5_DATA1_11) );
  DLH_X2 data_reg_10_ ( .G(n720), .D(ResultIn[2]), .Q(U5_DATA1_10) );
  DLH_X2 data_reg_9_ ( .G(n720), .D(ResultIn[1]), .Q(U5_DATA1_9) );
  DLH_X2 data_reg_8_ ( .G(n720), .D(ResultIn[0]), .Q(U5_DATA1_8) );
  DLH_X2 data_reg_7_ ( .G(n809), .D(ResultIn[7]), .Q(U5_DATA1_7) );
  DLH_X2 data_reg_6_ ( .G(n809), .D(ResultIn[6]), .Q(U5_DATA1_6) );
  DLH_X2 data_reg_5_ ( .G(n809), .D(ResultIn[5]), .Q(U5_DATA1_5) );
  DLH_X2 data_reg_4_ ( .G(n809), .D(ResultIn[4]), .Q(U5_DATA1_4) );
  DLH_X2 data_reg_3_ ( .G(n809), .D(ResultIn[3]), .Q(U5_DATA1_3) );
  DLH_X2 data_reg_2_ ( .G(n809), .D(ResultIn[2]), .Q(U5_DATA1_2) );
  DLH_X2 data_reg_1_ ( .G(n809), .D(ResultIn[1]), .Q(U5_DATA1_1) );
  DLH_X2 data_reg_0_ ( .G(n809), .D(ResultIn[0]), .Q(U5_DATA1_0) );
  DFF_X2 WriteAddress_reg_15_ ( .D(add_37_A_15_), .CK(clock), .Q(
        WriteAddress[15]) );
  DFF_X2 WriteAddress_reg_14_ ( .D(add_37_A_14_), .CK(clock), .Q(
        WriteAddress[14]) );
  DFF_X2 WriteAddress_reg_13_ ( .D(add_37_A_13_), .CK(clock), .Q(
        WriteAddress[13]) );
  DFF_X2 WriteAddress_reg_12_ ( .D(add_37_A_12_), .CK(clock), .Q(
        WriteAddress[12]) );
  DFF_X2 WriteAddress_reg_11_ ( .D(add_37_A_11_), .CK(clock), .Q(
        WriteAddress[11]) );
  DFF_X2 WriteAddress_reg_10_ ( .D(add_37_A_10_), .CK(clock), .Q(
        WriteAddress[10]) );
  DFF_X2 WriteAddress_reg_9_ ( .D(add_37_A_9_), .CK(clock), .Q(WriteAddress[9]) );
  DFF_X2 WriteAddress_reg_8_ ( .D(add_37_A_8_), .CK(clock), .Q(WriteAddress[8]) );
  DFF_X2 WriteAddress_reg_7_ ( .D(add_37_A_7_), .CK(clock), .Q(WriteAddress[7]) );
  DFF_X2 WriteAddress_reg_6_ ( .D(add_37_A_6_), .CK(clock), .Q(WriteAddress[6]) );
  DFF_X2 WriteAddress_reg_5_ ( .D(add_37_A_5_), .CK(clock), .Q(WriteAddress[5]) );
  DFFR_X2 next_WriteAddress_reg_5_ ( .D(n819), .CK(clock), .RN(n738), .Q(
        add_37_A_5_) );
  DFF_X2 WriteAddress_reg_4_ ( .D(add_37_A_4_), .CK(clock), .Q(WriteAddress[4]) );
  DFF_X2 WriteAddress_reg_3_ ( .D(add_37_A_3_), .CK(clock), .Q(WriteAddress[3]) );
  DFFR_X2 next_WriteAddress_reg_3_ ( .D(n821), .CK(clock), .RN(n738), .Q(
        add_37_A_3_) );
  DFF_X2 WriteAddress_reg_2_ ( .D(add_37_A_2_), .CK(clock), .Q(WriteAddress[2]) );
  DFF_X2 WriteAddress_reg_1_ ( .D(add_37_A_1_), .CK(clock), .Q(WriteAddress[1]) );
  DFFR_X2 next_WriteAddress_reg_1_ ( .D(n823), .CK(clock), .RN(n738), .Q(
        add_37_A_1_) );
  DFF_X2 WriteAddress_reg_0_ ( .D(add_37_A_0_), .CK(clock), .Q(WriteAddress[0]) );
  DFFR_X2 next_WriteAddress_reg_8_ ( .D(n816), .CK(clock), .RN(n737), .Q(
        add_37_A_8_), .QN(n772) );
  DFFR_X2 next_WriteAddress_reg_10_ ( .D(n814), .CK(clock), .RN(n738), .Q(
        add_37_A_10_), .QN(n781) );
  DFFR_X2 next_WriteAddress_reg_9_ ( .D(n815), .CK(clock), .RN(n738), .Q(
        add_37_A_9_) );
  DFFR_X2 next_WriteAddress_reg_7_ ( .D(n817), .CK(clock), .RN(n737), .Q(
        add_37_A_7_) );
  DFFR_X2 next_WriteAddress_reg_12_ ( .D(n812), .CK(clock), .RN(n737), .Q(
        add_37_A_12_), .QN(n790) );
  DFFR_X2 WriteEnable_reg ( .D(n733), .CK(clock), .RN(n738), .Q(WriteEnable)
         );
  DFFR_X2 next_WriteAddress_reg_6_ ( .D(n818), .CK(clock), .RN(n737), .Q(
        add_37_A_6_), .QN(n763) );
  DFFR_X2 next_WriteAddress_reg_11_ ( .D(n813), .CK(clock), .RN(n738), .Q(
        add_37_A_11_) );
  DFFR_X2 next_WriteAddress_reg_13_ ( .D(n811), .CK(clock), .RN(n737), .Q(
        add_37_A_13_), .QN(n798) );
  DFFR_X2 WriteBus_reg_9_ ( .D(n719), .CK(clock), .RN(reset_n), .Q(WriteBus[9]) );
  DFFR_X2 WriteBus_reg_8_ ( .D(n718), .CK(clock), .RN(n741), .Q(WriteBus[8])
         );
  DFFR_X2 WriteBus_reg_7_ ( .D(n717), .CK(clock), .RN(n738), .Q(WriteBus[7])
         );
  DFFR_X2 WriteBus_reg_6_ ( .D(n716), .CK(clock), .RN(n740), .Q(WriteBus[6])
         );
  DFFR_X2 WriteBus_reg_5_ ( .D(n715), .CK(clock), .RN(n741), .Q(WriteBus[5])
         );
  DFFR_X2 WriteBus_reg_4_ ( .D(n714), .CK(clock), .RN(n737), .Q(WriteBus[4])
         );
  DFFR_X2 WriteBus_reg_3_ ( .D(n713), .CK(clock), .RN(n740), .Q(WriteBus[3])
         );
  DFFR_X2 WriteBus_reg_2_ ( .D(n712), .CK(clock), .RN(n741), .Q(WriteBus[2])
         );
  DFFR_X2 WriteBus_reg_1_ ( .D(n711), .CK(clock), .RN(n738), .Q(WriteBus[1])
         );
  DFFR_X2 WriteBus_reg_25_ ( .D(n710), .CK(clock), .RN(n738), .Q(WriteBus[25])
         );
  DFFR_X2 WriteBus_reg_24_ ( .D(n709), .CK(clock), .RN(n740), .Q(WriteBus[24])
         );
  DFFR_X2 WriteBus_reg_23_ ( .D(n708), .CK(clock), .RN(n741), .Q(WriteBus[23])
         );
  DFFR_X2 WriteBus_reg_22_ ( .D(n707), .CK(clock), .RN(n737), .Q(WriteBus[22])
         );
  DFFR_X2 WriteBus_reg_21_ ( .D(n706), .CK(clock), .RN(n740), .Q(WriteBus[21])
         );
  DFFR_X2 WriteBus_reg_20_ ( .D(n705), .CK(clock), .RN(n741), .Q(WriteBus[20])
         );
  DFFR_X2 WriteBus_reg_19_ ( .D(n704), .CK(clock), .RN(n739), .Q(WriteBus[19])
         );
  DFFR_X2 WriteBus_reg_18_ ( .D(n703), .CK(clock), .RN(n740), .Q(WriteBus[18])
         );
  DFFR_X2 WriteBus_reg_17_ ( .D(n702), .CK(clock), .RN(n741), .Q(WriteBus[17])
         );
  DFFR_X2 WriteBus_reg_16_ ( .D(n701), .CK(clock), .RN(n738), .Q(WriteBus[16])
         );
  DFFR_X2 WriteBus_reg_15_ ( .D(n700), .CK(clock), .RN(n740), .Q(WriteBus[15])
         );
  DFFR_X2 WriteBus_reg_14_ ( .D(n699), .CK(clock), .RN(n741), .Q(WriteBus[14])
         );
  DFFR_X2 WriteBus_reg_13_ ( .D(n698), .CK(clock), .RN(n737), .Q(WriteBus[13])
         );
  DFFR_X2 WriteBus_reg_124_ ( .D(n697), .CK(clock), .RN(n737), .Q(
        WriteBus[124]) );
  DFFR_X2 WriteBus_reg_123_ ( .D(n696), .CK(clock), .RN(n738), .Q(
        WriteBus[123]) );
  DFFR_X2 WriteBus_reg_122_ ( .D(n695), .CK(clock), .RN(n737), .Q(
        WriteBus[122]) );
  DFFR_X2 WriteBus_reg_121_ ( .D(n694), .CK(clock), .RN(n738), .Q(
        WriteBus[121]) );
  DFFR_X2 WriteBus_reg_120_ ( .D(n693), .CK(clock), .RN(n737), .Q(
        WriteBus[120]) );
  DFFR_X2 WriteBus_reg_119_ ( .D(n692), .CK(clock), .RN(n738), .Q(
        WriteBus[119]) );
  DFFR_X2 WriteBus_reg_118_ ( .D(n691), .CK(clock), .RN(n737), .Q(
        WriteBus[118]) );
  DFFR_X2 WriteBus_reg_117_ ( .D(n690), .CK(clock), .RN(n738), .Q(
        WriteBus[117]) );
  DFFR_X2 WriteBus_reg_116_ ( .D(n689), .CK(clock), .RN(n738), .Q(
        WriteBus[116]) );
  DFFR_X2 WriteBus_reg_115_ ( .D(n688), .CK(clock), .RN(n737), .Q(
        WriteBus[115]) );
  DFFR_X2 WriteBus_reg_114_ ( .D(n687), .CK(clock), .RN(n738), .Q(
        WriteBus[114]) );
  DFFR_X2 WriteBus_reg_113_ ( .D(n686), .CK(clock), .RN(n737), .Q(
        WriteBus[113]) );
  DFFR_X2 WriteBus_reg_112_ ( .D(n685), .CK(clock), .RN(n738), .Q(
        WriteBus[112]) );
  DFFR_X2 WriteBus_reg_111_ ( .D(n684), .CK(clock), .RN(n737), .Q(
        WriteBus[111]) );
  DFFR_X2 WriteBus_reg_110_ ( .D(n683), .CK(clock), .RN(n738), .Q(
        WriteBus[110]) );
  DFFR_X2 WriteBus_reg_109_ ( .D(n682), .CK(clock), .RN(n737), .Q(
        WriteBus[109]) );
  DFFR_X2 WriteBus_reg_108_ ( .D(n681), .CK(clock), .RN(n738), .Q(
        WriteBus[108]) );
  DFFR_X2 WriteBus_reg_107_ ( .D(n680), .CK(clock), .RN(n737), .Q(
        WriteBus[107]) );
  DFFR_X2 WriteBus_reg_106_ ( .D(n679), .CK(clock), .RN(n739), .Q(
        WriteBus[106]) );
  DFFR_X2 WriteBus_reg_105_ ( .D(n678), .CK(clock), .RN(n739), .Q(
        WriteBus[105]) );
  DFFR_X2 WriteBus_reg_104_ ( .D(n677), .CK(clock), .RN(n739), .Q(
        WriteBus[104]) );
  DFFR_X2 WriteBus_reg_103_ ( .D(n676), .CK(clock), .RN(n739), .Q(
        WriteBus[103]) );
  DFFR_X2 WriteBus_reg_102_ ( .D(n675), .CK(clock), .RN(n739), .Q(
        WriteBus[102]) );
  DFFR_X2 WriteBus_reg_101_ ( .D(n674), .CK(clock), .RN(n739), .Q(
        WriteBus[101]) );
  DFFR_X2 WriteBus_reg_100_ ( .D(n673), .CK(clock), .RN(n739), .Q(
        WriteBus[100]) );
  DFFR_X2 WriteBus_reg_99_ ( .D(n672), .CK(clock), .RN(n739), .Q(WriteBus[99])
         );
  DFFR_X2 WriteBus_reg_98_ ( .D(n671), .CK(clock), .RN(n739), .Q(WriteBus[98])
         );
  DFFR_X2 WriteBus_reg_97_ ( .D(n670), .CK(clock), .RN(n739), .Q(WriteBus[97])
         );
  DFFR_X2 WriteBus_reg_96_ ( .D(n669), .CK(clock), .RN(n739), .Q(WriteBus[96])
         );
  DFFR_X2 WriteBus_reg_95_ ( .D(n668), .CK(clock), .RN(n739), .Q(WriteBus[95])
         );
  DFFR_X2 WriteBus_reg_94_ ( .D(n667), .CK(clock), .RN(n739), .Q(WriteBus[94])
         );
  DFFR_X2 WriteBus_reg_93_ ( .D(n666), .CK(clock), .RN(n739), .Q(WriteBus[93])
         );
  DFFR_X2 WriteBus_reg_92_ ( .D(n665), .CK(clock), .RN(n739), .Q(WriteBus[92])
         );
  DFFR_X2 WriteBus_reg_91_ ( .D(n664), .CK(clock), .RN(n739), .Q(WriteBus[91])
         );
  DFFR_X2 WriteBus_reg_90_ ( .D(n663), .CK(clock), .RN(n739), .Q(WriteBus[90])
         );
  DFFR_X2 WriteBus_reg_89_ ( .D(n662), .CK(clock), .RN(n739), .Q(WriteBus[89])
         );
  DFFR_X2 WriteBus_reg_88_ ( .D(n661), .CK(clock), .RN(n739), .Q(WriteBus[88])
         );
  DFFR_X2 WriteBus_reg_87_ ( .D(n660), .CK(clock), .RN(n740), .Q(WriteBus[87])
         );
  DFFR_X2 WriteBus_reg_86_ ( .D(n659), .CK(clock), .RN(n741), .Q(WriteBus[86])
         );
  DFFR_X2 WriteBus_reg_85_ ( .D(n658), .CK(clock), .RN(n737), .Q(WriteBus[85])
         );
  DFFR_X2 WriteBus_reg_84_ ( .D(n657), .CK(clock), .RN(n740), .Q(WriteBus[84])
         );
  DFFR_X2 WriteBus_reg_83_ ( .D(n656), .CK(clock), .RN(n741), .Q(WriteBus[83])
         );
  DFFR_X2 WriteBus_reg_82_ ( .D(n655), .CK(clock), .RN(n740), .Q(WriteBus[82])
         );
  DFFR_X2 WriteBus_reg_81_ ( .D(n654), .CK(clock), .RN(n740), .Q(WriteBus[81])
         );
  DFFR_X2 WriteBus_reg_80_ ( .D(n653), .CK(clock), .RN(n741), .Q(WriteBus[80])
         );
  DFFR_X2 WriteBus_reg_79_ ( .D(n652), .CK(clock), .RN(n738), .Q(WriteBus[79])
         );
  DFFR_X2 WriteBus_reg_78_ ( .D(n651), .CK(clock), .RN(n740), .Q(WriteBus[78])
         );
  DFFR_X2 WriteBus_reg_77_ ( .D(n650), .CK(clock), .RN(n741), .Q(WriteBus[77])
         );
  DFFR_X2 WriteBus_reg_76_ ( .D(n649), .CK(clock), .RN(n739), .Q(WriteBus[76])
         );
  DFFR_X2 WriteBus_reg_75_ ( .D(n648), .CK(clock), .RN(n740), .Q(WriteBus[75])
         );
  DFFR_X2 WriteBus_reg_74_ ( .D(n647), .CK(clock), .RN(n741), .Q(WriteBus[74])
         );
  DFFR_X2 WriteBus_reg_73_ ( .D(n646), .CK(clock), .RN(n737), .Q(WriteBus[73])
         );
  DFFR_X2 WriteBus_reg_72_ ( .D(n645), .CK(clock), .RN(n740), .Q(WriteBus[72])
         );
  DFFR_X2 WriteBus_reg_71_ ( .D(n644), .CK(clock), .RN(n741), .Q(WriteBus[71])
         );
  DFFR_X2 WriteBus_reg_70_ ( .D(n643), .CK(clock), .RN(n738), .Q(WriteBus[70])
         );
  DFFR_X2 WriteBus_reg_69_ ( .D(n642), .CK(clock), .RN(n740), .Q(WriteBus[69])
         );
  DFFR_X2 WriteBus_reg_68_ ( .D(n641), .CK(clock), .RN(n741), .Q(WriteBus[68])
         );
  DFFR_X2 WriteBus_reg_67_ ( .D(n640), .CK(clock), .RN(n739), .Q(WriteBus[67])
         );
  DFFR_X2 WriteBus_reg_66_ ( .D(n639), .CK(clock), .RN(n740), .Q(WriteBus[66])
         );
  DFFR_X2 WriteBus_reg_65_ ( .D(n638), .CK(clock), .RN(n741), .Q(WriteBus[65])
         );
  DFFR_X2 WriteBus_reg_64_ ( .D(n637), .CK(clock), .RN(n737), .Q(WriteBus[64])
         );
  DFFR_X2 WriteBus_reg_63_ ( .D(n636), .CK(clock), .RN(n740), .Q(WriteBus[63])
         );
  DFFR_X2 WriteBus_reg_62_ ( .D(n635), .CK(clock), .RN(n741), .Q(WriteBus[62])
         );
  DFFR_X2 WriteBus_reg_61_ ( .D(n634), .CK(clock), .RN(n739), .Q(WriteBus[61])
         );
  DFFR_X2 WriteBus_reg_60_ ( .D(n633), .CK(clock), .RN(n740), .Q(WriteBus[60])
         );
  DFFR_X2 WriteBus_reg_59_ ( .D(n632), .CK(clock), .RN(n741), .Q(WriteBus[59])
         );
  DFFR_X2 WriteBus_reg_58_ ( .D(n631), .CK(clock), .RN(n739), .Q(WriteBus[58])
         );
  DFFR_X2 WriteBus_reg_57_ ( .D(n630), .CK(clock), .RN(n740), .Q(WriteBus[57])
         );
  DFFR_X2 WriteBus_reg_56_ ( .D(n629), .CK(clock), .RN(n741), .Q(WriteBus[56])
         );
  DFFR_X2 WriteBus_reg_55_ ( .D(n628), .CK(clock), .RN(n738), .Q(WriteBus[55])
         );
  DFFR_X2 WriteBus_reg_54_ ( .D(n627), .CK(clock), .RN(n740), .Q(WriteBus[54])
         );
  DFFR_X2 WriteBus_reg_53_ ( .D(n626), .CK(clock), .RN(n741), .Q(WriteBus[53])
         );
  DFFR_X2 WriteBus_reg_52_ ( .D(n625), .CK(clock), .RN(n738), .Q(WriteBus[52])
         );
  DFFR_X2 WriteBus_reg_51_ ( .D(n624), .CK(clock), .RN(n740), .Q(WriteBus[51])
         );
  DFFR_X2 WriteBus_reg_50_ ( .D(n623), .CK(clock), .RN(n741), .Q(WriteBus[50])
         );
  DFFR_X2 WriteBus_reg_49_ ( .D(n622), .CK(clock), .RN(n739), .Q(WriteBus[49])
         );
  DFFR_X2 WriteBus_reg_48_ ( .D(n621), .CK(clock), .RN(n740), .Q(WriteBus[48])
         );
  DFFR_X2 WriteBus_reg_47_ ( .D(n620), .CK(clock), .RN(n741), .Q(WriteBus[47])
         );
  DFFR_X2 WriteBus_reg_46_ ( .D(n619), .CK(clock), .RN(n737), .Q(WriteBus[46])
         );
  DFFR_X2 WriteBus_reg_45_ ( .D(n618), .CK(clock), .RN(n740), .Q(WriteBus[45])
         );
  DFFR_X2 WriteBus_reg_44_ ( .D(n617), .CK(clock), .RN(n741), .Q(WriteBus[44])
         );
  DFFR_X2 WriteBus_reg_43_ ( .D(n616), .CK(clock), .RN(n738), .Q(WriteBus[43])
         );
  DFFR_X2 WriteBus_reg_42_ ( .D(n615), .CK(clock), .RN(n740), .Q(WriteBus[42])
         );
  DFFR_X2 WriteBus_reg_41_ ( .D(n614), .CK(clock), .RN(n741), .Q(WriteBus[41])
         );
  DFFR_X2 WriteBus_reg_40_ ( .D(n613), .CK(clock), .RN(n737), .Q(WriteBus[40])
         );
  DFFR_X2 WriteBus_reg_39_ ( .D(n612), .CK(clock), .RN(n740), .Q(WriteBus[39])
         );
  DFFR_X2 WriteBus_reg_38_ ( .D(n611), .CK(clock), .RN(n741), .Q(WriteBus[38])
         );
  DFFR_X2 WriteBus_reg_37_ ( .D(n610), .CK(clock), .RN(n739), .Q(WriteBus[37])
         );
  DFFR_X2 WriteBus_reg_36_ ( .D(n609), .CK(clock), .RN(n740), .Q(WriteBus[36])
         );
  DFFR_X2 WriteBus_reg_35_ ( .D(n608), .CK(clock), .RN(n741), .Q(WriteBus[35])
         );
  DFFR_X2 WriteBus_reg_34_ ( .D(n607), .CK(clock), .RN(n738), .Q(WriteBus[34])
         );
  DFFR_X2 WriteBus_reg_33_ ( .D(n606), .CK(clock), .RN(n740), .Q(WriteBus[33])
         );
  DFFR_X2 WriteBus_reg_32_ ( .D(n605), .CK(clock), .RN(n741), .Q(WriteBus[32])
         );
  DFFR_X2 WriteBus_reg_31_ ( .D(n604), .CK(clock), .RN(n737), .Q(WriteBus[31])
         );
  DFFR_X2 WriteBus_reg_30_ ( .D(n603), .CK(clock), .RN(n740), .Q(WriteBus[30])
         );
  DFFR_X2 WriteBus_reg_29_ ( .D(n602), .CK(clock), .RN(n741), .Q(WriteBus[29])
         );
  DFFR_X2 WriteBus_reg_28_ ( .D(n601), .CK(clock), .RN(n739), .Q(WriteBus[28])
         );
  DFFR_X2 WriteBus_reg_27_ ( .D(n600), .CK(clock), .RN(n740), .Q(WriteBus[27])
         );
  DFFR_X2 WriteBus_reg_26_ ( .D(n599), .CK(clock), .RN(n741), .Q(WriteBus[26])
         );
  DFFR_X2 WriteBus_reg_0_ ( .D(n598), .CK(clock), .RN(n741), .Q(WriteBus[0])
         );
  DFFR_X2 next_WriteAddress_reg_14_ ( .D(n810), .CK(clock), .RN(reset_n), .Q(
        add_37_A_14_) );
  DFFR_X2 next_WriteAddress_reg_15_ ( .D(n181), .CK(clock), .RN(reset_n), .Q(
        add_37_A_15_), .QN(n149) );
  DFFR_X2 WriteBus_reg_12_ ( .D(n597), .CK(clock), .RN(reset_n), .Q(
        WriteBus[12]) );
  DFFR_X2 WriteBus_reg_11_ ( .D(n596), .CK(clock), .RN(n739), .Q(WriteBus[11])
         );
  DFFR_X2 WriteBus_reg_10_ ( .D(n595), .CK(clock), .RN(n740), .Q(WriteBus[10])
         );
  DFFR_X2 WriteBus_reg_127_ ( .D(n594), .CK(clock), .RN(n737), .Q(
        WriteBus[127]) );
  DFFR_X2 WriteBus_reg_126_ ( .D(n593), .CK(clock), .RN(n738), .Q(
        WriteBus[126]) );
  DFFR_X2 WriteBus_reg_125_ ( .D(n592), .CK(clock), .RN(n737), .Q(
        WriteBus[125]) );
  DFFR_X1 next_WriteAddress_reg_0_ ( .D(n182), .CK(clock), .RN(n737), .Q(
        add_37_A_0_), .QN(n151) );
  DFFR_X1 next_WriteAddress_reg_4_ ( .D(n820), .CK(clock), .RN(n737), .Q(
        add_37_A_4_), .QN(n586) );
  DFFR_X1 next_WriteAddress_reg_2_ ( .D(n822), .CK(clock), .RN(n737), .Q(
        add_37_A_2_), .QN(n585) );
  AND2_X4 U3 ( .A1(n180), .A2(n148), .ZN(n578) );
  INV_X2 U4 ( .A(n801), .ZN(n733) );
  AND2_X4 U5 ( .A1(n731), .A2(n591), .ZN(n579) );
  AND2_X4 U6 ( .A1(n731), .A2(n590), .ZN(n580) );
  AND2_X4 U7 ( .A1(n730), .A2(n591), .ZN(n581) );
  AND2_X4 U8 ( .A1(n730), .A2(n590), .ZN(n582) );
  AND2_X4 U9 ( .A1(n732), .A2(n591), .ZN(n583) );
  AND2_X4 U10 ( .A1(n732), .A2(n590), .ZN(n584) );
  AND2_X4 U11 ( .A1(n729), .A2(n731), .ZN(n587) );
  AND2_X4 U12 ( .A1(n729), .A2(n730), .ZN(n588) );
  AND2_X4 U13 ( .A1(n729), .A2(n732), .ZN(n589) );
  AND2_X4 U14 ( .A1(sub_46_A_0_), .A2(n177), .ZN(n590) );
  AND2_X4 U15 ( .A1(n177), .A2(n148), .ZN(n591) );
  INV_X8 U16 ( .A(n742), .ZN(n741) );
  INV_X8 U17 ( .A(n742), .ZN(n740) );
  INV_X8 U18 ( .A(n742), .ZN(n739) );
  INV_X8 U19 ( .A(n742), .ZN(n738) );
  INV_X8 U20 ( .A(n742), .ZN(n737) );
  AND2_X1 U21 ( .A1(U5_DATA1_125), .A2(n734), .ZN(n592) );
  AND2_X1 U22 ( .A1(U5_DATA1_126), .A2(n733), .ZN(n593) );
  AND2_X1 U23 ( .A1(U5_DATA1_127), .A2(n734), .ZN(n594) );
  AND2_X1 U24 ( .A1(U5_DATA1_10), .A2(n734), .ZN(n595) );
  AND2_X1 U25 ( .A1(U5_DATA1_11), .A2(n734), .ZN(n596) );
  AND2_X1 U26 ( .A1(U5_DATA1_12), .A2(n734), .ZN(n597) );
  AND2_X1 U27 ( .A1(U5_DATA1_0), .A2(n735), .ZN(n598) );
  AND2_X1 U28 ( .A1(U5_DATA1_26), .A2(n734), .ZN(n599) );
  AND2_X1 U29 ( .A1(U5_DATA1_27), .A2(n734), .ZN(n600) );
  AND2_X1 U30 ( .A1(U5_DATA1_28), .A2(n735), .ZN(n601) );
  AND2_X1 U31 ( .A1(U5_DATA1_29), .A2(n733), .ZN(n602) );
  AND2_X1 U32 ( .A1(U5_DATA1_30), .A2(n734), .ZN(n603) );
  AND2_X1 U33 ( .A1(U5_DATA1_31), .A2(n733), .ZN(n604) );
  AND2_X1 U34 ( .A1(U5_DATA1_32), .A2(n735), .ZN(n605) );
  AND2_X1 U35 ( .A1(U5_DATA1_33), .A2(n734), .ZN(n606) );
  AND2_X1 U36 ( .A1(U5_DATA1_34), .A2(n734), .ZN(n607) );
  AND2_X1 U37 ( .A1(U5_DATA1_35), .A2(n733), .ZN(n608) );
  AND2_X1 U38 ( .A1(U5_DATA1_36), .A2(n735), .ZN(n609) );
  AND2_X1 U39 ( .A1(U5_DATA1_37), .A2(n734), .ZN(n610) );
  AND2_X1 U40 ( .A1(U5_DATA1_38), .A2(n733), .ZN(n611) );
  AND2_X1 U41 ( .A1(U5_DATA1_39), .A2(n734), .ZN(n612) );
  AND2_X1 U42 ( .A1(U5_DATA1_40), .A2(n735), .ZN(n613) );
  AND2_X1 U43 ( .A1(U5_DATA1_41), .A2(n734), .ZN(n614) );
  AND2_X1 U44 ( .A1(U5_DATA1_42), .A2(n734), .ZN(n615) );
  AND2_X1 U45 ( .A1(U5_DATA1_43), .A2(n733), .ZN(n616) );
  AND2_X1 U46 ( .A1(U5_DATA1_44), .A2(n735), .ZN(n617) );
  AND2_X1 U47 ( .A1(U5_DATA1_45), .A2(n734), .ZN(n618) );
  AND2_X1 U48 ( .A1(U5_DATA1_46), .A2(n734), .ZN(n619) );
  AND2_X1 U49 ( .A1(U5_DATA1_47), .A2(n734), .ZN(n620) );
  AND2_X1 U50 ( .A1(U5_DATA1_48), .A2(n735), .ZN(n621) );
  AND2_X1 U51 ( .A1(U5_DATA1_49), .A2(n733), .ZN(n622) );
  AND2_X1 U52 ( .A1(U5_DATA1_50), .A2(n734), .ZN(n623) );
  AND2_X1 U53 ( .A1(U5_DATA1_51), .A2(n735), .ZN(n624) );
  AND2_X1 U54 ( .A1(U5_DATA1_52), .A2(n734), .ZN(n625) );
  AND2_X1 U55 ( .A1(U5_DATA1_53), .A2(n734), .ZN(n626) );
  AND2_X1 U56 ( .A1(U5_DATA1_54), .A2(n734), .ZN(n627) );
  AND2_X1 U57 ( .A1(U5_DATA1_55), .A2(n735), .ZN(n628) );
  AND2_X1 U58 ( .A1(U5_DATA1_56), .A2(n734), .ZN(n629) );
  AND2_X1 U59 ( .A1(U5_DATA1_57), .A2(n734), .ZN(n630) );
  AND2_X1 U60 ( .A1(U5_DATA1_58), .A2(n734), .ZN(n631) );
  AND2_X1 U61 ( .A1(U5_DATA1_59), .A2(n735), .ZN(n632) );
  AND2_X1 U62 ( .A1(U5_DATA1_60), .A2(n734), .ZN(n633) );
  AND2_X1 U63 ( .A1(U5_DATA1_61), .A2(n733), .ZN(n634) );
  AND2_X1 U64 ( .A1(U5_DATA1_62), .A2(n733), .ZN(n635) );
  AND2_X1 U65 ( .A1(U5_DATA1_63), .A2(n735), .ZN(n636) );
  AND2_X1 U66 ( .A1(U5_DATA1_64), .A2(n734), .ZN(n637) );
  AND2_X1 U67 ( .A1(U5_DATA1_65), .A2(n735), .ZN(n638) );
  AND2_X1 U68 ( .A1(U5_DATA1_66), .A2(n735), .ZN(n639) );
  AND2_X1 U69 ( .A1(U5_DATA1_67), .A2(n735), .ZN(n640) );
  AND2_X1 U70 ( .A1(U5_DATA1_68), .A2(n735), .ZN(n641) );
  AND2_X1 U71 ( .A1(U5_DATA1_69), .A2(n735), .ZN(n642) );
  AND2_X1 U72 ( .A1(U5_DATA1_70), .A2(n735), .ZN(n643) );
  AND2_X1 U73 ( .A1(U5_DATA1_71), .A2(n735), .ZN(n644) );
  AND2_X1 U74 ( .A1(U5_DATA1_72), .A2(n735), .ZN(n645) );
  AND2_X1 U75 ( .A1(U5_DATA1_73), .A2(n735), .ZN(n646) );
  AND2_X1 U76 ( .A1(U5_DATA1_74), .A2(n735), .ZN(n647) );
  AND2_X1 U77 ( .A1(U5_DATA1_75), .A2(n735), .ZN(n648) );
  AND2_X1 U78 ( .A1(U5_DATA1_76), .A2(n735), .ZN(n649) );
  AND2_X1 U79 ( .A1(U5_DATA1_77), .A2(n734), .ZN(n650) );
  AND2_X1 U80 ( .A1(U5_DATA1_78), .A2(n733), .ZN(n651) );
  AND2_X1 U81 ( .A1(U5_DATA1_79), .A2(n734), .ZN(n652) );
  AND2_X1 U82 ( .A1(U5_DATA1_80), .A2(n733), .ZN(n653) );
  AND2_X1 U83 ( .A1(U5_DATA1_81), .A2(n734), .ZN(n654) );
  AND2_X1 U84 ( .A1(U5_DATA1_82), .A2(n734), .ZN(n655) );
  AND2_X1 U85 ( .A1(U5_DATA1_83), .A2(n734), .ZN(n656) );
  AND2_X1 U86 ( .A1(U5_DATA1_84), .A2(n734), .ZN(n657) );
  AND2_X1 U87 ( .A1(U5_DATA1_85), .A2(n734), .ZN(n658) );
  AND2_X1 U88 ( .A1(U5_DATA1_86), .A2(n733), .ZN(n659) );
  AND2_X1 U89 ( .A1(U5_DATA1_87), .A2(n735), .ZN(n660) );
  AND2_X1 U90 ( .A1(U5_DATA1_88), .A2(n734), .ZN(n661) );
  AND2_X1 U91 ( .A1(U5_DATA1_89), .A2(n734), .ZN(n662) );
  AND2_X1 U92 ( .A1(U5_DATA1_90), .A2(n735), .ZN(n663) );
  AND2_X1 U93 ( .A1(U5_DATA1_91), .A2(n733), .ZN(n664) );
  AND2_X1 U94 ( .A1(U5_DATA1_92), .A2(n735), .ZN(n665) );
  AND2_X1 U95 ( .A1(U5_DATA1_93), .A2(n735), .ZN(n666) );
  AND2_X1 U96 ( .A1(U5_DATA1_94), .A2(n734), .ZN(n667) );
  AND2_X1 U97 ( .A1(U5_DATA1_95), .A2(n735), .ZN(n668) );
  AND2_X1 U98 ( .A1(U5_DATA1_96), .A2(n734), .ZN(n669) );
  AND2_X1 U99 ( .A1(U5_DATA1_97), .A2(n734), .ZN(n670) );
  AND2_X1 U100 ( .A1(U5_DATA1_98), .A2(n735), .ZN(n671) );
  AND2_X1 U101 ( .A1(U5_DATA1_99), .A2(n734), .ZN(n672) );
  AND2_X1 U102 ( .A1(U5_DATA1_100), .A2(n734), .ZN(n673) );
  AND2_X1 U103 ( .A1(U5_DATA1_101), .A2(n735), .ZN(n674) );
  AND2_X1 U104 ( .A1(U5_DATA1_102), .A2(n735), .ZN(n675) );
  AND2_X1 U105 ( .A1(U5_DATA1_103), .A2(n734), .ZN(n676) );
  AND2_X1 U106 ( .A1(U5_DATA1_104), .A2(n734), .ZN(n677) );
  AND2_X1 U107 ( .A1(U5_DATA1_105), .A2(n734), .ZN(n678) );
  AND2_X1 U108 ( .A1(U5_DATA1_106), .A2(n733), .ZN(n679) );
  AND2_X1 U109 ( .A1(U5_DATA1_107), .A2(n734), .ZN(n680) );
  AND2_X1 U110 ( .A1(U5_DATA1_108), .A2(n734), .ZN(n681) );
  AND2_X1 U111 ( .A1(U5_DATA1_109), .A2(n734), .ZN(n682) );
  AND2_X1 U112 ( .A1(U5_DATA1_110), .A2(n734), .ZN(n683) );
  AND2_X1 U113 ( .A1(U5_DATA1_111), .A2(n733), .ZN(n684) );
  AND2_X1 U114 ( .A1(U5_DATA1_112), .A2(n734), .ZN(n685) );
  AND2_X1 U115 ( .A1(U5_DATA1_113), .A2(n734), .ZN(n686) );
  AND2_X1 U116 ( .A1(U5_DATA1_114), .A2(n734), .ZN(n687) );
  AND2_X1 U117 ( .A1(U5_DATA1_115), .A2(n734), .ZN(n688) );
  AND2_X1 U118 ( .A1(U5_DATA1_116), .A2(n735), .ZN(n689) );
  AND2_X1 U119 ( .A1(U5_DATA1_117), .A2(n734), .ZN(n690) );
  AND2_X1 U120 ( .A1(U5_DATA1_118), .A2(n734), .ZN(n691) );
  AND2_X1 U121 ( .A1(U5_DATA1_119), .A2(n734), .ZN(n692) );
  AND2_X1 U122 ( .A1(U5_DATA1_120), .A2(n735), .ZN(n693) );
  AND2_X1 U123 ( .A1(U5_DATA1_121), .A2(n734), .ZN(n694) );
  AND2_X1 U124 ( .A1(U5_DATA1_122), .A2(n735), .ZN(n695) );
  AND2_X1 U125 ( .A1(U5_DATA1_123), .A2(n733), .ZN(n696) );
  AND2_X1 U126 ( .A1(U5_DATA1_124), .A2(n735), .ZN(n697) );
  AND2_X1 U127 ( .A1(U5_DATA1_13), .A2(n735), .ZN(n698) );
  AND2_X1 U128 ( .A1(U5_DATA1_14), .A2(n734), .ZN(n699) );
  AND2_X1 U129 ( .A1(U5_DATA1_15), .A2(n735), .ZN(n700) );
  AND2_X1 U130 ( .A1(U5_DATA1_16), .A2(n735), .ZN(n701) );
  AND2_X1 U132 ( .A1(U5_DATA1_17), .A2(n733), .ZN(n702) );
  AND2_X1 U133 ( .A1(U5_DATA1_18), .A2(n734), .ZN(n703) );
  AND2_X1 U134 ( .A1(U5_DATA1_19), .A2(n735), .ZN(n704) );
  AND2_X1 U135 ( .A1(U5_DATA1_20), .A2(n734), .ZN(n705) );
  AND2_X1 U136 ( .A1(U5_DATA1_21), .A2(n734), .ZN(n706) );
  AND2_X1 U137 ( .A1(U5_DATA1_22), .A2(n735), .ZN(n707) );
  AND2_X1 U138 ( .A1(U5_DATA1_23), .A2(n734), .ZN(n708) );
  AND2_X1 U139 ( .A1(U5_DATA1_24), .A2(n735), .ZN(n709) );
  AND2_X1 U140 ( .A1(U5_DATA1_25), .A2(n735), .ZN(n710) );
  AND2_X1 U141 ( .A1(U5_DATA1_1), .A2(n734), .ZN(n711) );
  AND2_X1 U142 ( .A1(U5_DATA1_2), .A2(n734), .ZN(n712) );
  AND2_X1 U143 ( .A1(U5_DATA1_3), .A2(n734), .ZN(n713) );
  AND2_X1 U144 ( .A1(U5_DATA1_4), .A2(n734), .ZN(n714) );
  AND2_X1 U145 ( .A1(U5_DATA1_5), .A2(n734), .ZN(n715) );
  AND2_X1 U146 ( .A1(U5_DATA1_6), .A2(n734), .ZN(n716) );
  AND2_X1 U147 ( .A1(U5_DATA1_7), .A2(n734), .ZN(n717) );
  AND2_X1 U148 ( .A1(U5_DATA1_8), .A2(n734), .ZN(n718) );
  AND2_X1 U149 ( .A1(U5_DATA1_9), .A2(n734), .ZN(n719) );
  INV_X4 U150 ( .A(n736), .ZN(n735) );
  INV_X4 U151 ( .A(n733), .ZN(n736) );
  INV_X4 U152 ( .A(n801), .ZN(n734) );
  INV_X4 U153 ( .A(reset_n), .ZN(n742) );
  OAI21_X2 U154 ( .B1(n794), .B2(n801), .A(n155), .ZN(n797) );
  AND2_X1 U155 ( .A1(n727), .A2(n729), .ZN(n720) );
  AND2_X1 U156 ( .A1(n578), .A2(n731), .ZN(n721) );
  AND2_X1 U157 ( .A1(n578), .A2(n730), .ZN(n722) );
  AND2_X1 U158 ( .A1(n578), .A2(n732), .ZN(n723) );
  AND2_X1 U159 ( .A1(n727), .A2(n591), .ZN(n724) );
  AND2_X1 U160 ( .A1(n727), .A2(n590), .ZN(n725) );
  XOR2_X2 U162 ( .A(sub_46_A_4_), .B(n726), .Z(U4_DATA2_4) );
  NOR2_X1 U163 ( .A1(sub_46_A_3_), .A2(sub_46_carry_3_), .ZN(n726) );
  OAI21_X1 U164 ( .B1(n151), .B2(n155), .A(n744), .ZN(n182) );
  NOR2_X2 U165 ( .A1(sub_46_A_1_), .A2(sub_46_A_2_), .ZN(n727) );
  AND3_X2 U166 ( .A1(add_37_A_13_), .A2(n794), .A3(n734), .ZN(n728) );
  AND2_X1 U167 ( .A1(sub_46_A_0_), .A2(n180), .ZN(n729) );
  NOR2_X2 U168 ( .A1(n147), .A2(sub_46_A_1_), .ZN(n730) );
  AND2_X1 U169 ( .A1(sub_46_A_1_), .A2(n147), .ZN(n731) );
  AND2_X1 U170 ( .A1(sub_46_A_2_), .A2(sub_46_A_1_), .ZN(n732) );
  NAND2_X4 U171 ( .A1(StartIn), .A2(n809), .ZN(n801) );
  NAND2_X2 U173 ( .A1(n727), .A2(n578), .ZN(n743) );
  INV_X4 U174 ( .A(n743), .ZN(n809) );
  NAND2_X2 U175 ( .A1(StartIn), .A2(n801), .ZN(n155) );
  NAND2_X2 U176 ( .A1(n735), .A2(n151), .ZN(n744) );
  NOR2_X2 U178 ( .A1(n151), .A2(n801), .ZN(n745) );
  NAND2_X2 U179 ( .A1(n744), .A2(n155), .ZN(n747) );
  MUX2_X2 U180 ( .A(n745), .B(n747), .S(add_37_A_1_), .Z(n823) );
  NAND2_X2 U181 ( .A1(add_37_A_0_), .A2(n585), .ZN(n746) );
  MUX2_X2 U182 ( .A(n585), .B(n746), .S(add_37_A_1_), .Z(n749) );
  INV_X4 U183 ( .A(n747), .ZN(n748) );
  OAI22_X2 U184 ( .A1(n749), .A2(n801), .B1(n748), .B2(n585), .ZN(n822) );
  NAND3_X2 U185 ( .A1(add_37_A_1_), .A2(add_37_A_0_), .A3(add_37_A_2_), .ZN(
        n752) );
  NOR2_X2 U186 ( .A1(n752), .A2(n801), .ZN(n751) );
  NAND2_X2 U187 ( .A1(n735), .A2(n752), .ZN(n750) );
  NAND2_X2 U188 ( .A1(n750), .A2(n155), .ZN(n754) );
  MUX2_X2 U189 ( .A(n751), .B(n754), .S(add_37_A_3_), .Z(n821) );
  INV_X4 U190 ( .A(n752), .ZN(n757) );
  NAND2_X2 U191 ( .A1(n757), .A2(n586), .ZN(n753) );
  MUX2_X2 U192 ( .A(n586), .B(n753), .S(add_37_A_3_), .Z(n756) );
  INV_X4 U193 ( .A(n754), .ZN(n755) );
  OAI22_X2 U194 ( .A1(n756), .A2(n801), .B1(n755), .B2(n586), .ZN(n820) );
  NAND3_X2 U195 ( .A1(add_37_A_4_), .A2(add_37_A_3_), .A3(n757), .ZN(n760) );
  NOR2_X2 U199 ( .A1(n760), .A2(n801), .ZN(n759) );
  NAND2_X2 U200 ( .A1(n734), .A2(n760), .ZN(n758) );
  NAND2_X2 U201 ( .A1(n758), .A2(n155), .ZN(n762) );
  MUX2_X2 U202 ( .A(n759), .B(n762), .S(add_37_A_5_), .Z(n819) );
  INV_X4 U203 ( .A(n760), .ZN(n766) );
  NAND2_X2 U204 ( .A1(n766), .A2(n763), .ZN(n761) );
  MUX2_X2 U205 ( .A(n763), .B(n761), .S(add_37_A_5_), .Z(n765) );
  INV_X4 U206 ( .A(n762), .ZN(n764) );
  OAI22_X2 U207 ( .A1(n765), .A2(n801), .B1(n764), .B2(n763), .ZN(n818) );
  NAND3_X2 U208 ( .A1(add_37_A_6_), .A2(add_37_A_5_), .A3(n766), .ZN(n769) );
  NOR2_X2 U209 ( .A1(n769), .A2(n801), .ZN(n768) );
  NAND2_X2 U210 ( .A1(n735), .A2(n769), .ZN(n767) );
  NAND2_X2 U211 ( .A1(n767), .A2(n155), .ZN(n771) );
  MUX2_X2 U212 ( .A(n768), .B(n771), .S(add_37_A_7_), .Z(n817) );
  INV_X4 U213 ( .A(n769), .ZN(n775) );
  NAND2_X2 U214 ( .A1(n775), .A2(n772), .ZN(n770) );
  MUX2_X2 U215 ( .A(n772), .B(n770), .S(add_37_A_7_), .Z(n774) );
  INV_X4 U216 ( .A(n771), .ZN(n773) );
  OAI22_X2 U217 ( .A1(n774), .A2(n801), .B1(n773), .B2(n772), .ZN(n816) );
  NAND3_X2 U218 ( .A1(add_37_A_8_), .A2(add_37_A_7_), .A3(n775), .ZN(n778) );
  NOR2_X2 U219 ( .A1(n778), .A2(n801), .ZN(n777) );
  NAND2_X2 U220 ( .A1(n735), .A2(n778), .ZN(n776) );
  NAND2_X2 U221 ( .A1(n776), .A2(n155), .ZN(n780) );
  MUX2_X2 U222 ( .A(n777), .B(n780), .S(add_37_A_9_), .Z(n815) );
  INV_X4 U223 ( .A(n778), .ZN(n784) );
  NAND2_X2 U224 ( .A1(n784), .A2(n781), .ZN(n779) );
  MUX2_X2 U225 ( .A(n781), .B(n779), .S(add_37_A_9_), .Z(n783) );
  INV_X4 U226 ( .A(n780), .ZN(n782) );
  OAI22_X2 U227 ( .A1(n783), .A2(n801), .B1(n782), .B2(n781), .ZN(n814) );
  NAND3_X2 U228 ( .A1(add_37_A_10_), .A2(add_37_A_9_), .A3(n784), .ZN(n787) );
  NOR2_X2 U229 ( .A1(n787), .A2(n801), .ZN(n786) );
  NAND2_X2 U230 ( .A1(n734), .A2(n787), .ZN(n785) );
  NAND2_X2 U231 ( .A1(n785), .A2(n155), .ZN(n789) );
  MUX2_X2 U232 ( .A(n786), .B(n789), .S(add_37_A_11_), .Z(n813) );
  INV_X4 U233 ( .A(n787), .ZN(n793) );
  NAND2_X2 U234 ( .A1(n793), .A2(n790), .ZN(n788) );
  MUX2_X2 U235 ( .A(n790), .B(n788), .S(add_37_A_11_), .Z(n792) );
  INV_X4 U236 ( .A(n789), .ZN(n791) );
  OAI22_X2 U237 ( .A1(n792), .A2(n801), .B1(n791), .B2(n790), .ZN(n812) );
  NAND3_X2 U238 ( .A1(add_37_A_12_), .A2(add_37_A_11_), .A3(n793), .ZN(n796)
         );
  NOR2_X2 U239 ( .A1(n801), .A2(n796), .ZN(n795) );
  INV_X4 U240 ( .A(n796), .ZN(n794) );
  MUX2_X2 U241 ( .A(n795), .B(n797), .S(add_37_A_13_), .Z(n811) );
  INV_X4 U242 ( .A(n797), .ZN(n800) );
  NAND2_X2 U243 ( .A1(n733), .A2(n798), .ZN(n799) );
  NAND2_X2 U244 ( .A1(n800), .A2(n799), .ZN(n802) );
  MUX2_X2 U245 ( .A(n728), .B(n802), .S(add_37_A_14_), .Z(n810) );
  NAND3_X2 U246 ( .A1(output_base_offset), .A2(n801), .A3(n155), .ZN(n807) );
  NOR2_X2 U247 ( .A1(add_37_A_14_), .A2(n801), .ZN(n803) );
  NOR2_X2 U248 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X2 U249 ( .A1(add_37_A_14_), .A2(n728), .ZN(n804) );
  MUX2_X2 U250 ( .A(n805), .B(n804), .S(n149), .Z(n806) );
  NAND2_X2 U251 ( .A1(n807), .A2(n806), .ZN(n181) );
  INV_X4 U252 ( .A(n155), .ZN(n808) );
endmodule


module Output_top ( clock, reset_n, start, CdfMin, divisor, M2SP_ReadBus, 
        M2SP_ReadAddress, M3SP_ReadBus, M3SP_ReadAddress, WriteEnable, 
        Output_MEMBus, Output_MEMAddress, done, output_base_offset );
  input [19:0] CdfMin;
  input [19:0] divisor;
  input [127:0] M2SP_ReadBus;
  output [15:0] M2SP_ReadAddress;
  input [127:0] M3SP_ReadBus;
  output [15:0] M3SP_ReadAddress;
  output [127:0] Output_MEMBus;
  output [15:0] Output_MEMAddress;
  input clock, reset_n, start, output_base_offset;
  output WriteEnable, done;
  wire   start_to_stage_two, start_to_stage_three, start_to_stage_four,
         start_to_stage_five, n15, n16, n17, n18, n19, n20,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23;
  wire   [7:0] DataToStageTwo;
  wire   [19:0] DataToStageThree;
  wire   [27:0] DataToStageFour;
  wire   [7:0] result;
  assign M2SP_ReadAddress[14] = 1'b0;
  assign M2SP_ReadAddress[13] = 1'b0;
  assign M2SP_ReadAddress[12] = 1'b0;
  assign M2SP_ReadAddress[11] = 1'b0;
  assign M2SP_ReadAddress[10] = 1'b0;
  assign M2SP_ReadAddress[9] = 1'b0;
  assign M2SP_ReadAddress[8] = 1'b0;

  Output_Fetch_MEM stage1 ( .clock(clock), .reset_n(n19), .start(start), 
        .ReadBus(M3SP_ReadBus), .ReadAddress(M3SP_ReadAddress), .DataOut(
        DataToStageTwo), .StartOut(start_to_stage_two), .StoreAddress({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16}), .output_base_offset(n18), .done(done) );
  Output_Fetch_Cdf stage2 ( .clock(clock), .reset_n(n19), .ReadBus(
        M2SP_ReadBus), .ReadAddress({M2SP_ReadAddress[15], 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, M2SP_ReadAddress[7:0]}), .DataIn(
        DataToStageTwo), .DataOut(DataToStageThree), .StartIn(
        start_to_stage_two), .StartOut(start_to_stage_three), 
        .output_base_offset(n18) );
  Output_TopExpression stage3 ( .clock(clock), .reset_n(n19), .DataIn(
        DataToStageThree), .CdfMin({CdfMin[19:6], n16, CdfMin[4:0]}), 
        .StartIn(start_to_stage_three), .StartOut(start_to_stage_four), 
        .DataOut(DataToStageFour) );
  Output_Result stage4 ( .clock(clock), .reset_n(n19), .DataIn(DataToStageFour), .StartIn(start_to_stage_four), .Divisor(divisor), .StartOut(
        start_to_stage_five), .DataOut(result) );
  Output_Store stage5 ( .clock(clock), .reset_n(n19), .StartIn(
        start_to_stage_five), .ResultIn(result), .WriteBus(Output_MEMBus), 
        .WriteAddress(Output_MEMAddress), .WriteEnable(WriteEnable), 
        .output_base_offset(n18) );
  INV_X4 U16 ( .A(n15), .ZN(n16) );
  INV_X2 U17 ( .A(CdfMin[5]), .ZN(n15) );
  INV_X4 U18 ( .A(n17), .ZN(n18) );
  INV_X4 U19 ( .A(output_base_offset), .ZN(n17) );
  INV_X4 U20 ( .A(reset_n), .ZN(n20) );
  INV_X16 U1 ( .A(n20), .ZN(n19) );
endmodule


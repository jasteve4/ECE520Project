
module pipleline_stage_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(CO), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X4 U3 ( .A(B[0]), .ZN(n1) );
  INV_X4 U4 ( .A(A[0]), .ZN(n2) );
endmodule


module pipleline_stage_0 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n23;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;
  assign stage_out[7] = divided[6];
  assign stage_out[6] = divided[5];
  assign stage_out[5] = divided[4];
  assign stage_out[4] = divided[3];
  assign stage_out[3] = divided[2];
  assign stage_out[2] = divided[1];
  assign stage_out[1] = divided[0];

  pipleline_stage_0_DW01_add_0 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  XNOR2_X2 U4 ( .A(stage_result[20]), .B(divided[27]), .ZN(n23) );
  INV_X4 U5 ( .A(n23), .ZN(q) );
  MUX2_X1 U6 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9]) );
  MUX2_X1 U7 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8]) );
  MUX2_X1 U8 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27])
         );
  MUX2_X1 U9 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26])
         );
  MUX2_X1 U10 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X1 U11 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X1 U12 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X1 U13 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X1 U14 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X1 U15 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X1 U16 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X1 U17 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X1 U18 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X1 U19 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X1 U20 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X1 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X1 U22 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X1 U23 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X1 U24 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X1 U25 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
endmodule


module pipleline_stage_7_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(CO), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X4 U3 ( .A(B[0]), .ZN(n1) );
  INV_X4 U4 ( .A(A[0]), .ZN(n2) );
endmodule


module pipleline_stage_7 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n23;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;
  assign stage_out[7] = divided[6];
  assign stage_out[6] = divided[5];
  assign stage_out[5] = divided[4];
  assign stage_out[4] = divided[3];
  assign stage_out[3] = divided[2];
  assign stage_out[2] = divided[1];
  assign stage_out[1] = divided[0];

  pipleline_stage_7_DW01_add_0 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  XNOR2_X2 U4 ( .A(stage_result[20]), .B(divided[27]), .ZN(n23) );
  INV_X4 U5 ( .A(n23), .ZN(q) );
  MUX2_X1 U6 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9]) );
  MUX2_X1 U7 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8]) );
  MUX2_X1 U8 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27])
         );
  MUX2_X1 U9 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26])
         );
  MUX2_X1 U10 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X1 U11 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X1 U12 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X1 U13 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X1 U14 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X1 U15 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X1 U16 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X1 U17 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X1 U18 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X1 U19 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X1 U20 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X1 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X1 U22 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X1 U23 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X1 U24 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X1 U25 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
endmodule


module pipleline_stage_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(CO), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X4 U3 ( .A(B[0]), .ZN(n1) );
  INV_X4 U4 ( .A(A[0]), .ZN(n2) );
endmodule


module pipleline_stage_6 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n23;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;
  assign stage_out[7] = divided[6];
  assign stage_out[6] = divided[5];
  assign stage_out[5] = divided[4];
  assign stage_out[4] = divided[3];
  assign stage_out[3] = divided[2];
  assign stage_out[2] = divided[1];
  assign stage_out[1] = divided[0];

  pipleline_stage_6_DW01_add_0 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  XNOR2_X2 U4 ( .A(stage_result[20]), .B(divided[27]), .ZN(n23) );
  INV_X4 U5 ( .A(n23), .ZN(q) );
  MUX2_X1 U6 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9]) );
  MUX2_X1 U7 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8]) );
  MUX2_X1 U8 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27])
         );
  MUX2_X1 U9 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26])
         );
  MUX2_X1 U10 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X1 U11 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X1 U12 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X1 U13 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X1 U14 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X1 U15 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X1 U16 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X1 U17 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X1 U18 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X1 U19 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X1 U20 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X1 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X1 U22 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X1 U23 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X1 U24 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X1 U25 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
endmodule


module pipleline_stage_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(CO), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X4 U3 ( .A(B[0]), .ZN(n1) );
  INV_X4 U4 ( .A(A[0]), .ZN(n2) );
endmodule


module pipleline_stage_5 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n23;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;
  assign stage_out[7] = divided[6];
  assign stage_out[6] = divided[5];
  assign stage_out[5] = divided[4];
  assign stage_out[4] = divided[3];
  assign stage_out[3] = divided[2];
  assign stage_out[2] = divided[1];
  assign stage_out[1] = divided[0];

  pipleline_stage_5_DW01_add_0 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  XNOR2_X2 U4 ( .A(stage_result[20]), .B(divided[27]), .ZN(n23) );
  INV_X4 U5 ( .A(n23), .ZN(q) );
  MUX2_X1 U6 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9]) );
  MUX2_X1 U7 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8]) );
  MUX2_X1 U8 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27])
         );
  MUX2_X1 U9 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26])
         );
  MUX2_X1 U10 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X1 U11 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X1 U12 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X1 U13 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X1 U14 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X1 U15 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X1 U16 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X1 U17 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X1 U18 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X1 U19 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X1 U20 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X1 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X1 U22 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X1 U23 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X1 U24 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X1 U25 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
endmodule


module pipleline_stage_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(CO), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X4 U3 ( .A(B[0]), .ZN(n1) );
  INV_X4 U4 ( .A(A[0]), .ZN(n2) );
endmodule


module pipleline_stage_4 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n23;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;
  assign stage_out[7] = divided[6];
  assign stage_out[6] = divided[5];
  assign stage_out[5] = divided[4];
  assign stage_out[4] = divided[3];
  assign stage_out[3] = divided[2];
  assign stage_out[2] = divided[1];
  assign stage_out[1] = divided[0];

  pipleline_stage_4_DW01_add_0 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  XNOR2_X2 U4 ( .A(stage_result[20]), .B(divided[27]), .ZN(n23) );
  INV_X4 U5 ( .A(n23), .ZN(q) );
  MUX2_X1 U6 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9]) );
  MUX2_X1 U7 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8]) );
  MUX2_X1 U8 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27])
         );
  MUX2_X1 U9 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26])
         );
  MUX2_X1 U10 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X1 U11 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X1 U12 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X1 U13 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X1 U14 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X1 U15 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X1 U16 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X1 U17 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X1 U18 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X1 U19 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X1 U20 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X1 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X1 U22 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X1 U23 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X1 U24 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X1 U25 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
endmodule


module pipleline_stage_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(CO), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X4 U3 ( .A(B[0]), .ZN(n1) );
  INV_X4 U4 ( .A(A[0]), .ZN(n2) );
endmodule


module pipleline_stage_3 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n23;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;
  assign stage_out[7] = divided[6];
  assign stage_out[6] = divided[5];
  assign stage_out[5] = divided[4];
  assign stage_out[4] = divided[3];
  assign stage_out[3] = divided[2];
  assign stage_out[2] = divided[1];
  assign stage_out[1] = divided[0];

  pipleline_stage_3_DW01_add_0 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  XNOR2_X2 U4 ( .A(stage_result[20]), .B(divided[27]), .ZN(n23) );
  INV_X4 U5 ( .A(n23), .ZN(q) );
  MUX2_X1 U6 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9]) );
  MUX2_X1 U7 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8]) );
  MUX2_X1 U8 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27])
         );
  MUX2_X1 U9 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26])
         );
  MUX2_X1 U10 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X1 U11 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X1 U12 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X1 U13 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X1 U14 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X1 U15 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X1 U16 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X1 U17 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X1 U18 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X1 U19 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X1 U20 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X1 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X1 U22 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X1 U23 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X1 U24 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X1 U25 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
endmodule


module pipleline_stage_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(CO), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X4 U3 ( .A(B[0]), .ZN(n1) );
  INV_X4 U4 ( .A(A[0]), .ZN(n2) );
endmodule


module pipleline_stage_2 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n23;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;
  assign stage_out[7] = divided[6];
  assign stage_out[6] = divided[5];
  assign stage_out[5] = divided[4];
  assign stage_out[4] = divided[3];
  assign stage_out[3] = divided[2];
  assign stage_out[2] = divided[1];
  assign stage_out[1] = divided[0];

  pipleline_stage_2_DW01_add_0 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  XNOR2_X2 U4 ( .A(stage_result[20]), .B(divided[27]), .ZN(n23) );
  INV_X4 U5 ( .A(n23), .ZN(q) );
  MUX2_X1 U6 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9]) );
  MUX2_X1 U7 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8]) );
  MUX2_X1 U8 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27])
         );
  MUX2_X1 U9 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26])
         );
  MUX2_X1 U10 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X1 U11 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X1 U12 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X1 U13 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X1 U14 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X1 U15 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X1 U16 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X1 U17 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X1 U18 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X1 U19 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X1 U20 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X1 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X1 U22 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X1 U23 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X1 U24 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X1 U25 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
endmodule


module pipleline_stage_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [19:1] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(CO), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X4 U3 ( .A(B[0]), .ZN(n1) );
  INV_X4 U4 ( .A(A[0]), .ZN(n2) );
endmodule


module pipleline_stage_1 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n23;
  wire   [20:0] stage_result;
  assign stage_out[0] = 1'b0;
  assign stage_out[7] = divided[6];
  assign stage_out[6] = divided[5];
  assign stage_out[5] = divided[4];
  assign stage_out[4] = divided[3];
  assign stage_out[3] = divided[2];
  assign stage_out[2] = divided[1];
  assign stage_out[1] = divided[0];

  pipleline_stage_1_DW01_add_0 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  XNOR2_X2 U4 ( .A(stage_result[20]), .B(divided[27]), .ZN(n23) );
  INV_X4 U5 ( .A(n23), .ZN(q) );
  MUX2_X1 U6 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9]) );
  MUX2_X1 U7 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8]) );
  MUX2_X1 U8 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27])
         );
  MUX2_X1 U9 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26])
         );
  MUX2_X1 U10 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X1 U11 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X1 U12 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X1 U13 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X1 U14 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X1 U15 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X1 U16 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X1 U17 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X1 U18 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X1 U19 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X1 U20 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X1 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X1 U22 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X1 U23 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X1 U24 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X1 U25 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
endmodule


module pipeline_divider ( clock, reset_n, start, divided, divisor, q, StartOut
 );
  input [27:0] divided;
  input [19:0] divisor;
  output [7:0] q;
  input clock, reset_n, start;
  output StartOut;
  wire   q_bit7, StartOut0, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, N44, N65, q_bit6, StartOut1, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, q_bit5, StartOut2, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, q_bit4, StartOut3, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, q_bit3, StartOut4, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, q_bit2, StartOut5, N278, N279, N280, N281, N282, N283,
         N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294,
         N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305,
         N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316,
         N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327,
         N328, N329, N330, q_bit1, N333, N334, N335, N336, N337, N338, N339,
         N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350,
         N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361,
         N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372,
         N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
         N384, N385, N386, q_bit0, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35;
  wire   [27:1] stage0_result;
  wire   [27:0] pipe0_result;
  wire   [19:0] pipe0_divisor_n;
  wire   [27:1] stage1_result;
  wire   [27:0] pipe1_result;
  wire   [19:0] pipe1_divisor_n;
  wire   [27:1] stage2_result;
  wire   [27:0] pipe2_result;
  wire   [19:0] pipe2_divisor_n;
  wire   [27:1] stage3_result;
  wire   [27:0] pipe3_result;
  wire   [19:0] pipe3_divisor_n;
  wire   [27:1] stage4_result;
  wire   [27:0] pipe4_result;
  wire   [19:0] pipe4_divisor_n;
  wire   [27:1] stage5_result;
  wire   [27:0] pipe5_result;
  wire   [19:0] pipe5_divisor_n;
  wire   [27:1] stage6_result;
  wire   [27:0] pipe6_result;
  wire   [19:0] pipe6_divisor_n;

  pipleline_stage_0 stage0 ( .divided(divided), .divisor({n226, n227, n228, 
        n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
        n241, n242, n243, n244, n245}), .q(q_bit7), .stage_out({stage0_result, 
        SYNOPSYS_UNCONNECTED_1}) );
  pipleline_stage_7 stage1 ( .divided({pipe0_result[27:1], 1'b0}), .divisor(
        pipe0_divisor_n), .q(q_bit6), .stage_out({stage1_result, 
        SYNOPSYS_UNCONNECTED_2}) );
  pipleline_stage_6 stage2 ( .divided({pipe1_result[27:1], 1'b0}), .divisor(
        pipe1_divisor_n), .q(q_bit5), .stage_out({stage2_result, 
        SYNOPSYS_UNCONNECTED_3}) );
  pipleline_stage_5 stage3 ( .divided({pipe2_result[27:1], 1'b0}), .divisor(
        pipe2_divisor_n), .q(q_bit4), .stage_out({stage3_result, 
        SYNOPSYS_UNCONNECTED_4}) );
  pipleline_stage_4 stage4 ( .divided({pipe3_result[27:1], 1'b0}), .divisor(
        pipe3_divisor_n), .q(q_bit3), .stage_out({stage4_result, 
        SYNOPSYS_UNCONNECTED_5}) );
  pipleline_stage_3 stage5 ( .divided({pipe4_result[27:1], 1'b0}), .divisor(
        pipe4_divisor_n), .q(q_bit2), .stage_out({stage5_result, 
        SYNOPSYS_UNCONNECTED_6}) );
  pipleline_stage_2 stage6 ( .divided({pipe5_result[27:1], 1'b0}), .divisor(
        pipe5_divisor_n), .q(q_bit1), .stage_out({stage6_result, 
        SYNOPSYS_UNCONNECTED_7}) );
  pipleline_stage_1 stage7 ( .divided({pipe6_result[27:1], 1'b0}), .divisor(
        pipe6_divisor_n), .q(q_bit0), .stage_out({SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35}) );
  SDFFR_X2 pipe0_divisor_n_reg_19_ ( .D(1'b0), .SI(start), .SE(n226), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[19]), .QN(n210) );
  SDFFR_X2 pipe0_divisor_n_reg_18_ ( .D(1'b0), .SI(start), .SE(n227), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[18]), .QN(n211) );
  SDFFR_X2 pipe0_divisor_n_reg_17_ ( .D(1'b0), .SI(start), .SE(n228), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[17]), .QN(n212) );
  SDFFR_X2 pipe0_divisor_n_reg_16_ ( .D(1'b0), .SI(start), .SE(n229), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[16]), .QN(n213) );
  SDFFR_X2 pipe0_divisor_n_reg_15_ ( .D(1'b0), .SI(start), .SE(n230), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[15]), .QN(n214) );
  SDFFR_X2 pipe0_divisor_n_reg_14_ ( .D(1'b0), .SI(start), .SE(n231), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[14]), .QN(n215) );
  SDFFR_X2 pipe0_divisor_n_reg_13_ ( .D(1'b0), .SI(start), .SE(n232), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[13]), .QN(n216) );
  SDFFR_X2 pipe0_divisor_n_reg_12_ ( .D(1'b0), .SI(start), .SE(n233), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[12]), .QN(n217) );
  SDFFR_X2 pipe0_divisor_n_reg_11_ ( .D(1'b0), .SI(start), .SE(n234), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[11]), .QN(n218) );
  SDFFR_X2 pipe0_divisor_n_reg_10_ ( .D(1'b0), .SI(start), .SE(n235), .CK(
        clock), .RN(reset_n), .Q(pipe0_divisor_n[10]), .QN(n219) );
  SDFFR_X2 pipe0_divisor_n_reg_9_ ( .D(1'b0), .SI(start), .SE(n236), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[9]), .QN(n220) );
  SDFFR_X2 pipe0_divisor_n_reg_8_ ( .D(1'b0), .SI(start), .SE(n237), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[8]), .QN(n221) );
  SDFFR_X2 pipe0_divisor_n_reg_7_ ( .D(1'b0), .SI(start), .SE(n238), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[7]), .QN(n222) );
  SDFFR_X2 pipe0_divisor_n_reg_6_ ( .D(1'b0), .SI(start), .SE(n239), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[6]), .QN(n223) );
  SDFFR_X2 pipe0_divisor_n_reg_5_ ( .D(1'b0), .SI(start), .SE(n240), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[5]), .QN(n225) );
  SDFFR_X2 pipe0_divisor_n_reg_4_ ( .D(1'b0), .SI(start), .SE(n241), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[4]), .QN(n79) );
  SDFFR_X2 pipe0_divisor_n_reg_3_ ( .D(1'b0), .SI(start), .SE(n242), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[3]), .QN(n80) );
  SDFFR_X2 pipe0_divisor_n_reg_2_ ( .D(1'b0), .SI(start), .SE(n243), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[2]), .QN(n81) );
  SDFFR_X2 pipe0_divisor_n_reg_1_ ( .D(1'b0), .SI(start), .SE(n244), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[1]), .QN(n82) );
  SDFFR_X2 pipe0_divisor_n_reg_0_ ( .D(1'b0), .SI(start), .SE(n245), .CK(clock), .RN(reset_n), .Q(pipe0_divisor_n[0]), .QN(n83) );
  DFFR_X1 pipe0_q_reg_0_ ( .D(N65), .CK(clock), .RN(reset_n), .QN(n209) );
  DFFR_X1 pipe0_result_reg_27_ ( .D(N44), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[27]) );
  DFFR_X1 pipe0_result_reg_26_ ( .D(N43), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[26]) );
  DFFR_X1 pipe0_result_reg_25_ ( .D(N42), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[25]) );
  DFFR_X1 pipe0_result_reg_24_ ( .D(N41), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[24]) );
  DFFR_X1 pipe0_result_reg_23_ ( .D(N40), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[23]) );
  DFFR_X1 pipe0_result_reg_22_ ( .D(N39), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[22]) );
  DFFR_X1 pipe0_result_reg_21_ ( .D(N38), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[21]) );
  DFFR_X1 pipe0_result_reg_20_ ( .D(N37), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[20]) );
  DFFR_X1 pipe0_result_reg_19_ ( .D(N36), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[19]) );
  DFFR_X1 pipe0_result_reg_18_ ( .D(N35), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[18]) );
  DFFR_X1 pipe0_result_reg_17_ ( .D(N34), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[17]) );
  DFFR_X1 pipe0_result_reg_16_ ( .D(N33), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[16]) );
  DFFR_X1 pipe0_result_reg_15_ ( .D(N32), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[15]) );
  DFFR_X1 pipe0_result_reg_14_ ( .D(N31), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[14]) );
  DFFR_X1 pipe0_result_reg_13_ ( .D(N30), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[13]) );
  DFFR_X1 pipe0_result_reg_12_ ( .D(N29), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[12]) );
  DFFR_X1 pipe0_result_reg_11_ ( .D(N28), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[11]) );
  DFFR_X1 pipe0_result_reg_10_ ( .D(N27), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[10]) );
  DFFR_X1 pipe0_result_reg_9_ ( .D(N26), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[9]) );
  DFFR_X1 pipe0_result_reg_8_ ( .D(N25), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[8]) );
  DFFR_X1 pipe0_result_reg_7_ ( .D(N24), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[7]) );
  DFFR_X1 pipe0_result_reg_6_ ( .D(N23), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[6]) );
  DFFR_X1 pipe0_result_reg_5_ ( .D(N22), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[5]) );
  DFFR_X1 pipe0_result_reg_4_ ( .D(N21), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[4]) );
  DFFR_X1 pipe0_result_reg_3_ ( .D(N20), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[3]) );
  DFFR_X1 pipe0_result_reg_2_ ( .D(N19), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[2]) );
  DFFR_X1 pipe0_result_reg_1_ ( .D(N18), .CK(clock), .RN(reset_n), .Q(
        pipe0_result[1]) );
  DFFR_X1 pipe1_divisor_n_reg_19_ ( .D(N114), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[19]), .QN(n188) );
  DFFR_X1 pipe1_divisor_n_reg_18_ ( .D(N113), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[18]), .QN(n189) );
  DFFR_X1 pipe1_divisor_n_reg_17_ ( .D(N112), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[17]), .QN(n190) );
  DFFR_X1 pipe1_divisor_n_reg_16_ ( .D(N111), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[16]), .QN(n191) );
  DFFR_X1 pipe1_divisor_n_reg_15_ ( .D(N110), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[15]), .QN(n192) );
  DFFR_X1 pipe1_divisor_n_reg_14_ ( .D(N109), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[14]), .QN(n193) );
  DFFR_X1 pipe1_divisor_n_reg_13_ ( .D(N108), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[13]), .QN(n194) );
  DFFR_X1 pipe1_divisor_n_reg_12_ ( .D(N107), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[12]), .QN(n195) );
  DFFR_X1 pipe1_divisor_n_reg_11_ ( .D(N106), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[11]), .QN(n196) );
  DFFR_X1 pipe1_divisor_n_reg_10_ ( .D(N105), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[10]), .QN(n197) );
  DFFR_X1 pipe1_divisor_n_reg_9_ ( .D(N104), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[9]), .QN(n198) );
  DFFR_X1 pipe1_divisor_n_reg_8_ ( .D(N103), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[8]), .QN(n199) );
  DFFR_X1 pipe1_divisor_n_reg_7_ ( .D(N102), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[7]), .QN(n200) );
  DFFR_X1 pipe1_divisor_n_reg_6_ ( .D(N101), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[6]), .QN(n201) );
  DFFR_X1 pipe1_divisor_n_reg_5_ ( .D(N100), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[5]), .QN(n202) );
  DFFR_X1 pipe1_divisor_n_reg_4_ ( .D(N99), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[4]), .QN(n203) );
  DFFR_X1 pipe1_divisor_n_reg_3_ ( .D(N98), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[3]), .QN(n204) );
  DFFR_X1 pipe1_divisor_n_reg_2_ ( .D(N97), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[2]), .QN(n205) );
  DFFR_X1 pipe1_divisor_n_reg_1_ ( .D(N96), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[1]), .QN(n206) );
  DFFR_X1 pipe1_divisor_n_reg_0_ ( .D(N95), .CK(clock), .RN(reset_n), .Q(
        pipe1_divisor_n[0]), .QN(n207) );
  DFFR_X1 pipe1_q_reg_1_ ( .D(N116), .CK(clock), .RN(reset_n), .QN(n186) );
  DFFR_X1 pipe1_q_reg_0_ ( .D(N115), .CK(clock), .RN(reset_n), .QN(n187) );
  DFFR_X1 pipe1_result_reg_27_ ( .D(N94), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[27]) );
  DFFR_X1 pipe1_result_reg_26_ ( .D(N93), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[26]) );
  DFFR_X1 pipe1_result_reg_25_ ( .D(N92), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[25]) );
  DFFR_X1 pipe1_result_reg_24_ ( .D(N91), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[24]) );
  DFFR_X1 pipe1_result_reg_23_ ( .D(N90), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[23]) );
  DFFR_X1 pipe1_result_reg_22_ ( .D(N89), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[22]) );
  DFFR_X1 pipe1_result_reg_21_ ( .D(N88), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[21]) );
  DFFR_X1 pipe1_result_reg_20_ ( .D(N87), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[20]) );
  DFFR_X1 pipe1_result_reg_19_ ( .D(N86), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[19]) );
  DFFR_X1 pipe1_result_reg_18_ ( .D(N85), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[18]) );
  DFFR_X1 pipe1_result_reg_17_ ( .D(N84), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[17]) );
  DFFR_X1 pipe1_result_reg_16_ ( .D(N83), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[16]) );
  DFFR_X1 pipe1_result_reg_15_ ( .D(N82), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[15]) );
  DFFR_X1 pipe1_result_reg_14_ ( .D(N81), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[14]) );
  DFFR_X1 pipe1_result_reg_13_ ( .D(N80), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[13]) );
  DFFR_X1 pipe1_result_reg_12_ ( .D(N79), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[12]) );
  DFFR_X1 pipe1_result_reg_11_ ( .D(N78), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[11]) );
  DFFR_X1 pipe1_result_reg_10_ ( .D(N77), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[10]) );
  DFFR_X1 pipe1_result_reg_9_ ( .D(N76), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[9]) );
  DFFR_X1 pipe1_result_reg_8_ ( .D(N75), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[8]) );
  DFFR_X1 pipe1_result_reg_7_ ( .D(N74), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[7]) );
  DFFR_X1 pipe1_result_reg_6_ ( .D(N73), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[6]) );
  DFFR_X1 pipe1_result_reg_5_ ( .D(N72), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[5]) );
  DFFR_X1 pipe1_result_reg_4_ ( .D(N71), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[4]) );
  DFFR_X1 pipe1_result_reg_3_ ( .D(N70), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[3]) );
  DFFR_X1 pipe1_result_reg_2_ ( .D(N69), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[2]) );
  DFFR_X1 pipe1_result_reg_1_ ( .D(N68), .CK(clock), .RN(reset_n), .Q(
        pipe1_result[1]) );
  DFFR_X1 pipe2_divisor_n_reg_19_ ( .D(N165), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[19]), .QN(n165) );
  DFFR_X1 pipe2_divisor_n_reg_18_ ( .D(N164), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[18]), .QN(n166) );
  DFFR_X1 pipe2_divisor_n_reg_17_ ( .D(N163), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[17]), .QN(n167) );
  DFFR_X1 pipe2_divisor_n_reg_16_ ( .D(N162), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[16]), .QN(n168) );
  DFFR_X1 pipe2_divisor_n_reg_15_ ( .D(N161), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[15]), .QN(n169) );
  DFFR_X1 pipe2_divisor_n_reg_14_ ( .D(N160), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[14]), .QN(n170) );
  DFFR_X1 pipe2_divisor_n_reg_13_ ( .D(N159), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[13]), .QN(n171) );
  DFFR_X1 pipe2_divisor_n_reg_12_ ( .D(N158), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[12]), .QN(n172) );
  DFFR_X1 pipe2_divisor_n_reg_11_ ( .D(N157), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[11]), .QN(n173) );
  DFFR_X1 pipe2_divisor_n_reg_10_ ( .D(N156), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[10]), .QN(n174) );
  DFFR_X1 pipe2_divisor_n_reg_9_ ( .D(N155), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[9]), .QN(n175) );
  DFFR_X1 pipe2_divisor_n_reg_8_ ( .D(N154), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[8]), .QN(n176) );
  DFFR_X1 pipe2_divisor_n_reg_7_ ( .D(N153), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[7]), .QN(n177) );
  DFFR_X1 pipe2_divisor_n_reg_6_ ( .D(N152), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[6]), .QN(n178) );
  DFFR_X1 pipe2_divisor_n_reg_5_ ( .D(N151), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[5]), .QN(n179) );
  DFFR_X1 pipe2_divisor_n_reg_4_ ( .D(N150), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[4]), .QN(n180) );
  DFFR_X1 pipe2_divisor_n_reg_3_ ( .D(N149), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[3]), .QN(n181) );
  DFFR_X1 pipe2_divisor_n_reg_2_ ( .D(N148), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[2]), .QN(n182) );
  DFFR_X1 pipe2_divisor_n_reg_1_ ( .D(N147), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[1]), .QN(n183) );
  DFFR_X1 pipe2_divisor_n_reg_0_ ( .D(N146), .CK(clock), .RN(reset_n), .Q(
        pipe2_divisor_n[0]), .QN(n184) );
  DFFR_X1 pipe2_q_reg_2_ ( .D(N168), .CK(clock), .RN(reset_n), .QN(n162) );
  DFFR_X1 pipe2_q_reg_1_ ( .D(N167), .CK(clock), .RN(reset_n), .QN(n163) );
  DFFR_X1 pipe2_q_reg_0_ ( .D(N166), .CK(clock), .RN(reset_n), .QN(n164) );
  DFFR_X1 pipe2_result_reg_27_ ( .D(N145), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[27]) );
  DFFR_X1 pipe2_result_reg_26_ ( .D(N144), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[26]) );
  DFFR_X1 pipe2_result_reg_25_ ( .D(N143), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[25]) );
  DFFR_X1 pipe2_result_reg_24_ ( .D(N142), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[24]) );
  DFFR_X1 pipe2_result_reg_23_ ( .D(N141), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[23]) );
  DFFR_X1 pipe2_result_reg_22_ ( .D(N140), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[22]) );
  DFFR_X1 pipe2_result_reg_21_ ( .D(N139), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[21]) );
  DFFR_X1 pipe2_result_reg_20_ ( .D(N138), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[20]) );
  DFFR_X1 pipe2_result_reg_19_ ( .D(N137), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[19]) );
  DFFR_X1 pipe2_result_reg_18_ ( .D(N136), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[18]) );
  DFFR_X1 pipe2_result_reg_17_ ( .D(N135), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[17]) );
  DFFR_X1 pipe2_result_reg_16_ ( .D(N134), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[16]) );
  DFFR_X1 pipe2_result_reg_15_ ( .D(N133), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[15]) );
  DFFR_X1 pipe2_result_reg_14_ ( .D(N132), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[14]) );
  DFFR_X1 pipe2_result_reg_13_ ( .D(N131), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[13]) );
  DFFR_X1 pipe2_result_reg_12_ ( .D(N130), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[12]) );
  DFFR_X1 pipe2_result_reg_11_ ( .D(N129), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[11]) );
  DFFR_X1 pipe2_result_reg_10_ ( .D(N128), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[10]) );
  DFFR_X1 pipe2_result_reg_9_ ( .D(N127), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[9]) );
  DFFR_X1 pipe2_result_reg_8_ ( .D(N126), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[8]) );
  DFFR_X1 pipe2_result_reg_7_ ( .D(N125), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[7]) );
  DFFR_X1 pipe2_result_reg_6_ ( .D(N124), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[6]) );
  DFFR_X1 pipe2_result_reg_5_ ( .D(N123), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[5]) );
  DFFR_X1 pipe2_result_reg_4_ ( .D(N122), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[4]) );
  DFFR_X1 pipe2_result_reg_3_ ( .D(N121), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[3]) );
  DFFR_X1 pipe2_result_reg_2_ ( .D(N120), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[2]) );
  DFFR_X1 pipe2_result_reg_1_ ( .D(N119), .CK(clock), .RN(reset_n), .Q(
        pipe2_result[1]) );
  DFFR_X1 pipe3_divisor_n_reg_19_ ( .D(N217), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[19]), .QN(n141) );
  DFFR_X1 pipe3_divisor_n_reg_18_ ( .D(N216), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[18]), .QN(n142) );
  DFFR_X1 pipe3_divisor_n_reg_17_ ( .D(N215), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[17]), .QN(n143) );
  DFFR_X1 pipe3_divisor_n_reg_16_ ( .D(N214), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[16]), .QN(n144) );
  DFFR_X1 pipe3_divisor_n_reg_15_ ( .D(N213), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[15]), .QN(n145) );
  DFFR_X1 pipe3_divisor_n_reg_14_ ( .D(N212), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[14]), .QN(n146) );
  DFFR_X1 pipe3_divisor_n_reg_13_ ( .D(N211), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[13]), .QN(n147) );
  DFFR_X1 pipe3_divisor_n_reg_12_ ( .D(N210), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[12]), .QN(n148) );
  DFFR_X1 pipe3_divisor_n_reg_11_ ( .D(N209), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[11]), .QN(n149) );
  DFFR_X1 pipe3_divisor_n_reg_10_ ( .D(N208), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[10]), .QN(n150) );
  DFFR_X1 pipe3_divisor_n_reg_9_ ( .D(N207), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[9]), .QN(n151) );
  DFFR_X1 pipe3_divisor_n_reg_8_ ( .D(N206), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[8]), .QN(n152) );
  DFFR_X1 pipe3_divisor_n_reg_7_ ( .D(N205), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[7]), .QN(n153) );
  DFFR_X1 pipe3_divisor_n_reg_6_ ( .D(N204), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[6]), .QN(n154) );
  DFFR_X1 pipe3_divisor_n_reg_5_ ( .D(N203), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[5]), .QN(n155) );
  DFFR_X1 pipe3_divisor_n_reg_4_ ( .D(N202), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[4]), .QN(n156) );
  DFFR_X1 pipe3_divisor_n_reg_3_ ( .D(N201), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[3]), .QN(n157) );
  DFFR_X1 pipe3_divisor_n_reg_2_ ( .D(N200), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[2]), .QN(n158) );
  DFFR_X1 pipe3_divisor_n_reg_1_ ( .D(N199), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[1]), .QN(n159) );
  DFFR_X1 pipe3_divisor_n_reg_0_ ( .D(N198), .CK(clock), .RN(reset_n), .Q(
        pipe3_divisor_n[0]), .QN(n160) );
  DFFR_X1 pipe3_q_reg_3_ ( .D(N221), .CK(clock), .RN(reset_n), .QN(n137) );
  DFFR_X1 pipe3_q_reg_2_ ( .D(N220), .CK(clock), .RN(reset_n), .QN(n138) );
  DFFR_X1 pipe3_q_reg_1_ ( .D(N219), .CK(clock), .RN(reset_n), .QN(n139) );
  DFFR_X1 pipe3_q_reg_0_ ( .D(N218), .CK(clock), .RN(reset_n), .QN(n140) );
  DFFR_X1 pipe3_result_reg_27_ ( .D(N197), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[27]) );
  DFFR_X1 pipe3_result_reg_26_ ( .D(N196), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[26]) );
  DFFR_X1 pipe3_result_reg_25_ ( .D(N195), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[25]) );
  DFFR_X1 pipe3_result_reg_24_ ( .D(N194), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[24]) );
  DFFR_X1 pipe3_result_reg_23_ ( .D(N193), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[23]) );
  DFFR_X1 pipe3_result_reg_22_ ( .D(N192), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[22]) );
  DFFR_X1 pipe3_result_reg_21_ ( .D(N191), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[21]) );
  DFFR_X1 pipe3_result_reg_20_ ( .D(N190), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[20]) );
  DFFR_X1 pipe3_result_reg_19_ ( .D(N189), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[19]) );
  DFFR_X1 pipe3_result_reg_18_ ( .D(N188), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[18]) );
  DFFR_X1 pipe3_result_reg_17_ ( .D(N187), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[17]) );
  DFFR_X1 pipe3_result_reg_16_ ( .D(N186), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[16]) );
  DFFR_X1 pipe3_result_reg_15_ ( .D(N185), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[15]) );
  DFFR_X1 pipe3_result_reg_14_ ( .D(N184), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[14]) );
  DFFR_X1 pipe3_result_reg_13_ ( .D(N183), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[13]) );
  DFFR_X1 pipe3_result_reg_12_ ( .D(N182), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[12]) );
  DFFR_X1 pipe3_result_reg_11_ ( .D(N181), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[11]) );
  DFFR_X1 pipe3_result_reg_10_ ( .D(N180), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[10]) );
  DFFR_X1 pipe3_result_reg_9_ ( .D(N179), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[9]) );
  DFFR_X1 pipe3_result_reg_8_ ( .D(N178), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[8]) );
  DFFR_X1 pipe3_result_reg_7_ ( .D(N177), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[7]) );
  DFFR_X1 pipe3_result_reg_6_ ( .D(N176), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[6]) );
  DFFR_X1 pipe3_result_reg_5_ ( .D(N175), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[5]) );
  DFFR_X1 pipe3_result_reg_4_ ( .D(N174), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[4]) );
  DFFR_X1 pipe3_result_reg_3_ ( .D(N173), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[3]) );
  DFFR_X1 pipe3_result_reg_2_ ( .D(N172), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[2]) );
  DFFR_X1 pipe3_result_reg_1_ ( .D(N171), .CK(clock), .RN(reset_n), .Q(
        pipe3_result[1]) );
  DFFR_X1 pipe4_divisor_n_reg_19_ ( .D(N270), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[19]), .QN(n116) );
  DFFR_X1 pipe4_divisor_n_reg_18_ ( .D(N269), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[18]), .QN(n117) );
  DFFR_X1 pipe4_divisor_n_reg_17_ ( .D(N268), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[17]), .QN(n118) );
  DFFR_X1 pipe4_divisor_n_reg_16_ ( .D(N267), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[16]), .QN(n119) );
  DFFR_X1 pipe4_divisor_n_reg_15_ ( .D(N266), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[15]), .QN(n120) );
  DFFR_X1 pipe4_divisor_n_reg_14_ ( .D(N265), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[14]), .QN(n121) );
  DFFR_X1 pipe4_divisor_n_reg_13_ ( .D(N264), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[13]), .QN(n122) );
  DFFR_X1 pipe4_divisor_n_reg_12_ ( .D(N263), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[12]), .QN(n123) );
  DFFR_X1 pipe4_divisor_n_reg_11_ ( .D(N262), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[11]), .QN(n124) );
  DFFR_X1 pipe4_divisor_n_reg_10_ ( .D(N261), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[10]), .QN(n125) );
  DFFR_X1 pipe4_divisor_n_reg_9_ ( .D(N260), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[9]), .QN(n126) );
  DFFR_X1 pipe4_divisor_n_reg_8_ ( .D(N259), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[8]), .QN(n127) );
  DFFR_X1 pipe4_divisor_n_reg_7_ ( .D(N258), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[7]), .QN(n128) );
  DFFR_X1 pipe4_divisor_n_reg_6_ ( .D(N257), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[6]), .QN(n129) );
  DFFR_X1 pipe4_divisor_n_reg_5_ ( .D(N256), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[5]), .QN(n130) );
  DFFR_X1 pipe4_divisor_n_reg_4_ ( .D(N255), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[4]), .QN(n131) );
  DFFR_X1 pipe4_divisor_n_reg_3_ ( .D(N254), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[3]), .QN(n132) );
  DFFR_X1 pipe4_divisor_n_reg_2_ ( .D(N253), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[2]), .QN(n133) );
  DFFR_X1 pipe4_divisor_n_reg_1_ ( .D(N252), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[1]), .QN(n134) );
  DFFR_X1 pipe4_divisor_n_reg_0_ ( .D(N251), .CK(clock), .RN(reset_n), .Q(
        pipe4_divisor_n[0]), .QN(n135) );
  DFFR_X1 pipe4_q_reg_4_ ( .D(N275), .CK(clock), .RN(reset_n), .QN(n111) );
  DFFR_X1 pipe4_q_reg_3_ ( .D(N274), .CK(clock), .RN(reset_n), .QN(n112) );
  DFFR_X1 pipe4_q_reg_2_ ( .D(N273), .CK(clock), .RN(reset_n), .QN(n113) );
  DFFR_X1 pipe4_q_reg_1_ ( .D(N272), .CK(clock), .RN(reset_n), .QN(n114) );
  DFFR_X1 pipe4_q_reg_0_ ( .D(N271), .CK(clock), .RN(reset_n), .QN(n115) );
  DFFR_X1 pipe4_result_reg_27_ ( .D(N250), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[27]) );
  DFFR_X1 pipe4_result_reg_26_ ( .D(N249), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[26]) );
  DFFR_X1 pipe4_result_reg_25_ ( .D(N248), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[25]) );
  DFFR_X1 pipe4_result_reg_24_ ( .D(N247), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[24]) );
  DFFR_X1 pipe4_result_reg_23_ ( .D(N246), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[23]) );
  DFFR_X1 pipe4_result_reg_22_ ( .D(N245), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[22]) );
  DFFR_X1 pipe4_result_reg_21_ ( .D(N244), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[21]) );
  DFFR_X1 pipe4_result_reg_20_ ( .D(N243), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[20]) );
  DFFR_X1 pipe4_result_reg_19_ ( .D(N242), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[19]) );
  DFFR_X1 pipe4_result_reg_18_ ( .D(N241), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[18]) );
  DFFR_X1 pipe4_result_reg_17_ ( .D(N240), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[17]) );
  DFFR_X1 pipe4_result_reg_16_ ( .D(N239), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[16]) );
  DFFR_X1 pipe4_result_reg_15_ ( .D(N238), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[15]) );
  DFFR_X1 pipe4_result_reg_14_ ( .D(N237), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[14]) );
  DFFR_X1 pipe4_result_reg_13_ ( .D(N236), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[13]) );
  DFFR_X1 pipe4_result_reg_12_ ( .D(N235), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[12]) );
  DFFR_X1 pipe4_result_reg_11_ ( .D(N234), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[11]) );
  DFFR_X1 pipe4_result_reg_10_ ( .D(N233), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[10]) );
  DFFR_X1 pipe4_result_reg_9_ ( .D(N232), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[9]) );
  DFFR_X1 pipe4_result_reg_8_ ( .D(N231), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[8]) );
  DFFR_X1 pipe4_result_reg_7_ ( .D(N230), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[7]) );
  DFFR_X1 pipe4_result_reg_6_ ( .D(N229), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[6]) );
  DFFR_X1 pipe4_result_reg_5_ ( .D(N228), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[5]) );
  DFFR_X1 pipe4_result_reg_4_ ( .D(N227), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[4]) );
  DFFR_X1 pipe4_result_reg_3_ ( .D(N226), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[3]) );
  DFFR_X1 pipe4_result_reg_2_ ( .D(N225), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[2]) );
  DFFR_X1 pipe4_result_reg_1_ ( .D(N224), .CK(clock), .RN(reset_n), .Q(
        pipe4_result[1]) );
  DFFR_X1 pipe5_divisor_n_reg_19_ ( .D(N324), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[19]), .QN(n90) );
  DFFR_X1 pipe5_divisor_n_reg_18_ ( .D(N323), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[18]), .QN(n91) );
  DFFR_X1 pipe5_divisor_n_reg_17_ ( .D(N322), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[17]), .QN(n92) );
  DFFR_X1 pipe5_divisor_n_reg_16_ ( .D(N321), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[16]), .QN(n93) );
  DFFR_X1 pipe5_divisor_n_reg_15_ ( .D(N320), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[15]), .QN(n94) );
  DFFR_X1 pipe5_divisor_n_reg_14_ ( .D(N319), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[14]), .QN(n95) );
  DFFR_X1 pipe5_divisor_n_reg_13_ ( .D(N318), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[13]), .QN(n96) );
  DFFR_X1 pipe5_divisor_n_reg_12_ ( .D(N317), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[12]), .QN(n97) );
  DFFR_X1 pipe5_divisor_n_reg_11_ ( .D(N316), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[11]), .QN(n98) );
  DFFR_X1 pipe5_divisor_n_reg_10_ ( .D(N315), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[10]), .QN(n99) );
  DFFR_X1 pipe5_divisor_n_reg_9_ ( .D(N314), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[9]), .QN(n100) );
  DFFR_X1 pipe5_divisor_n_reg_8_ ( .D(N313), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[8]), .QN(n101) );
  DFFR_X1 pipe5_divisor_n_reg_7_ ( .D(N312), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[7]), .QN(n102) );
  DFFR_X1 pipe5_divisor_n_reg_6_ ( .D(N311), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[6]), .QN(n103) );
  DFFR_X1 pipe5_divisor_n_reg_5_ ( .D(N310), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[5]), .QN(n104) );
  DFFR_X1 pipe5_divisor_n_reg_4_ ( .D(N309), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[4]), .QN(n105) );
  DFFR_X1 pipe5_divisor_n_reg_3_ ( .D(N308), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[3]), .QN(n106) );
  DFFR_X1 pipe5_divisor_n_reg_2_ ( .D(N307), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[2]), .QN(n107) );
  DFFR_X1 pipe5_divisor_n_reg_1_ ( .D(N306), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[1]), .QN(n108) );
  DFFR_X1 pipe5_divisor_n_reg_0_ ( .D(N305), .CK(clock), .RN(reset_n), .Q(
        pipe5_divisor_n[0]), .QN(n109) );
  DFFR_X1 pipe5_q_reg_5_ ( .D(N330), .CK(clock), .RN(reset_n), .QN(n84) );
  DFFR_X1 pipe5_q_reg_4_ ( .D(N329), .CK(clock), .RN(reset_n), .QN(n85) );
  DFFR_X1 pipe5_q_reg_3_ ( .D(N328), .CK(clock), .RN(reset_n), .QN(n86) );
  DFFR_X1 pipe5_q_reg_2_ ( .D(N327), .CK(clock), .RN(reset_n), .QN(n87) );
  DFFR_X1 pipe5_q_reg_1_ ( .D(N326), .CK(clock), .RN(reset_n), .QN(n88) );
  DFFR_X1 pipe5_q_reg_0_ ( .D(N325), .CK(clock), .RN(reset_n), .QN(n89) );
  DFFR_X1 pipe5_result_reg_27_ ( .D(N304), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[27]) );
  DFFR_X1 pipe5_result_reg_26_ ( .D(N303), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[26]) );
  DFFR_X1 pipe5_result_reg_25_ ( .D(N302), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[25]) );
  DFFR_X1 pipe5_result_reg_24_ ( .D(N301), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[24]) );
  DFFR_X1 pipe5_result_reg_23_ ( .D(N300), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[23]) );
  DFFR_X1 pipe5_result_reg_22_ ( .D(N299), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[22]) );
  DFFR_X1 pipe5_result_reg_21_ ( .D(N298), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[21]) );
  DFFR_X1 pipe5_result_reg_20_ ( .D(N297), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[20]) );
  DFFR_X1 pipe5_result_reg_19_ ( .D(N296), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[19]) );
  DFFR_X1 pipe5_result_reg_18_ ( .D(N295), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[18]) );
  DFFR_X1 pipe5_result_reg_17_ ( .D(N294), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[17]) );
  DFFR_X1 pipe5_result_reg_16_ ( .D(N293), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[16]) );
  DFFR_X1 pipe5_result_reg_15_ ( .D(N292), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[15]) );
  DFFR_X1 pipe5_result_reg_14_ ( .D(N291), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[14]) );
  DFFR_X1 pipe5_result_reg_13_ ( .D(N290), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[13]) );
  DFFR_X1 pipe5_result_reg_12_ ( .D(N289), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[12]) );
  DFFR_X1 pipe5_result_reg_11_ ( .D(N288), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[11]) );
  DFFR_X1 pipe5_result_reg_10_ ( .D(N287), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[10]) );
  DFFR_X1 pipe5_result_reg_9_ ( .D(N286), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[9]) );
  DFFR_X1 pipe5_result_reg_8_ ( .D(N285), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[8]) );
  DFFR_X1 pipe5_result_reg_7_ ( .D(N284), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[7]) );
  DFFR_X1 pipe5_result_reg_6_ ( .D(N283), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[6]) );
  DFFR_X1 pipe5_result_reg_5_ ( .D(N282), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[5]) );
  DFFR_X1 pipe5_result_reg_4_ ( .D(N281), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[4]) );
  DFFR_X1 pipe5_result_reg_3_ ( .D(N280), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[3]) );
  DFFR_X1 pipe5_result_reg_2_ ( .D(N279), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[2]) );
  DFFR_X1 pipe5_result_reg_1_ ( .D(N278), .CK(clock), .RN(reset_n), .Q(
        pipe5_result[1]) );
  DFFR_X1 pipe6_divisor_n_reg_19_ ( .D(N379), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[19]) );
  DFFR_X1 pipe6_divisor_n_reg_18_ ( .D(N378), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[18]), .QN(n67) );
  DFFR_X1 pipe6_divisor_n_reg_17_ ( .D(N377), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[17]), .QN(n66) );
  DFFR_X1 pipe6_divisor_n_reg_16_ ( .D(N376), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[16]), .QN(n68) );
  DFFR_X1 pipe6_divisor_n_reg_15_ ( .D(N375), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[15]) );
  DFFR_X1 pipe6_divisor_n_reg_14_ ( .D(N374), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[14]) );
  DFFR_X1 pipe6_divisor_n_reg_13_ ( .D(N373), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[13]), .QN(n70) );
  DFFR_X1 pipe6_divisor_n_reg_12_ ( .D(N372), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[12]), .QN(n69) );
  DFFR_X1 pipe6_divisor_n_reg_11_ ( .D(N371), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[11]), .QN(n71) );
  DFFR_X1 pipe6_divisor_n_reg_10_ ( .D(N370), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[10]) );
  DFFR_X1 pipe6_divisor_n_reg_9_ ( .D(N369), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[9]), .QN(n61) );
  DFFR_X1 pipe6_divisor_n_reg_8_ ( .D(N368), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[8]), .QN(n60) );
  DFFR_X1 pipe6_divisor_n_reg_7_ ( .D(N367), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[7]), .QN(n62) );
  DFFR_X1 pipe6_divisor_n_reg_6_ ( .D(N366), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[6]) );
  DFFR_X1 pipe6_divisor_n_reg_5_ ( .D(N365), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[5]) );
  DFFR_X1 pipe6_divisor_n_reg_4_ ( .D(N364), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[4]), .QN(n64) );
  DFFR_X1 pipe6_divisor_n_reg_3_ ( .D(N363), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[3]), .QN(n63) );
  DFFR_X1 pipe6_divisor_n_reg_2_ ( .D(N362), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[2]), .QN(n65) );
  DFFR_X1 pipe6_divisor_n_reg_1_ ( .D(N361), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[1]) );
  DFFR_X1 pipe6_divisor_n_reg_0_ ( .D(N360), .CK(clock), .RN(reset_n), .Q(
        pipe6_divisor_n[0]) );
  DFFR_X1 pipe6_q_reg_6_ ( .D(N386), .CK(clock), .RN(reset_n), .QN(n72) );
  DFFR_X1 pipe6_q_reg_5_ ( .D(N385), .CK(clock), .RN(reset_n), .QN(n73) );
  DFFR_X1 pipe6_q_reg_4_ ( .D(N384), .CK(clock), .RN(reset_n), .QN(n74) );
  DFFR_X1 pipe6_q_reg_3_ ( .D(N383), .CK(clock), .RN(reset_n), .QN(n75) );
  DFFR_X1 pipe6_q_reg_2_ ( .D(N382), .CK(clock), .RN(reset_n), .QN(n76) );
  DFFR_X1 pipe6_q_reg_1_ ( .D(N381), .CK(clock), .RN(reset_n), .QN(n77) );
  DFFR_X1 pipe6_q_reg_0_ ( .D(N380), .CK(clock), .RN(reset_n), .QN(n78) );
  DFFR_X1 StartOut_reg ( .D(StartOut5), .CK(clock), .RN(reset_n), .Q(StartOut)
         );
  DFFR_X1 pipe6_result_reg_27_ ( .D(N359), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[27]) );
  DFFR_X1 pipe6_result_reg_26_ ( .D(N358), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[26]) );
  DFFR_X1 pipe6_result_reg_25_ ( .D(N357), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[25]) );
  DFFR_X1 pipe6_result_reg_24_ ( .D(N356), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[24]) );
  DFFR_X1 pipe6_result_reg_23_ ( .D(N355), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[23]) );
  DFFR_X1 pipe6_result_reg_22_ ( .D(N354), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[22]) );
  DFFR_X1 pipe6_result_reg_21_ ( .D(N353), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[21]) );
  DFFR_X1 pipe6_result_reg_20_ ( .D(N352), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[20]) );
  DFFR_X1 pipe6_result_reg_19_ ( .D(N351), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[19]) );
  DFFR_X1 pipe6_result_reg_18_ ( .D(N350), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[18]) );
  DFFR_X1 pipe6_result_reg_17_ ( .D(N349), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[17]) );
  DFFR_X1 pipe6_result_reg_16_ ( .D(N348), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[16]) );
  DFFR_X1 pipe6_result_reg_15_ ( .D(N347), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[15]) );
  DFFR_X1 pipe6_result_reg_14_ ( .D(N346), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[14]) );
  DFFR_X1 pipe6_result_reg_13_ ( .D(N345), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[13]) );
  DFFR_X1 pipe6_result_reg_12_ ( .D(N344), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[12]) );
  DFFR_X1 pipe6_result_reg_11_ ( .D(N343), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[11]) );
  DFFR_X1 pipe6_result_reg_10_ ( .D(N342), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[10]) );
  DFFR_X1 pipe6_result_reg_9_ ( .D(N341), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[9]) );
  DFFR_X1 pipe6_result_reg_8_ ( .D(N340), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[8]) );
  DFFR_X1 pipe6_result_reg_7_ ( .D(N339), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[7]) );
  DFFR_X1 pipe6_result_reg_6_ ( .D(N338), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[6]) );
  DFFR_X1 pipe6_result_reg_5_ ( .D(N337), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[5]) );
  DFFR_X1 pipe6_result_reg_4_ ( .D(N336), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[4]) );
  DFFR_X1 pipe6_result_reg_3_ ( .D(N335), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[3]) );
  DFFR_X1 pipe6_result_reg_2_ ( .D(N334), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[2]) );
  DFFR_X1 pipe6_result_reg_1_ ( .D(N333), .CK(clock), .RN(reset_n), .Q(
        pipe6_result[1]) );
  DFFR_X2 StartOut0_reg ( .D(start), .CK(clock), .RN(reset_n), .Q(StartOut0), 
        .QN(n224) );
  DFFR_X2 StartOut1_reg ( .D(StartOut0), .CK(clock), .RN(reset_n), .Q(
        StartOut1), .QN(n208) );
  DFFR_X2 StartOut2_reg ( .D(StartOut1), .CK(clock), .RN(reset_n), .Q(
        StartOut2), .QN(n185) );
  DFFR_X2 StartOut3_reg ( .D(StartOut2), .CK(clock), .RN(reset_n), .Q(
        StartOut3), .QN(n161) );
  DFFR_X2 StartOut4_reg ( .D(StartOut3), .CK(clock), .RN(reset_n), .Q(
        StartOut4), .QN(n136) );
  DFFR_X2 StartOut5_reg ( .D(StartOut4), .CK(clock), .RN(reset_n), .Q(
        StartOut5), .QN(n110) );
  NOR2_X1 U411 ( .A1(n50), .A2(n72), .ZN(q[7]) );
  NOR2_X1 U412 ( .A1(n50), .A2(n73), .ZN(q[6]) );
  NOR2_X1 U413 ( .A1(n50), .A2(n74), .ZN(q[5]) );
  NOR2_X1 U414 ( .A1(n50), .A2(n75), .ZN(q[4]) );
  NOR2_X1 U415 ( .A1(n50), .A2(n76), .ZN(q[3]) );
  NOR2_X1 U416 ( .A1(n50), .A2(n77), .ZN(q[2]) );
  NOR2_X1 U417 ( .A1(n50), .A2(n78), .ZN(q[1]) );
  INV_X1 U418 ( .A(n51), .ZN(n50) );
  AND2_X1 U419 ( .A1(q_bit0), .A2(n51), .ZN(q[0]) );
  NAND4_X1 U420 ( .A1(n52), .A2(n53), .A3(n54), .A4(n55), .ZN(n51) );
  NOR3_X1 U421 ( .A1(n56), .A2(pipe6_divisor_n[6]), .A3(pipe6_divisor_n[5]), 
        .ZN(n55) );
  NAND3_X1 U422 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n56) );
  NOR3_X1 U423 ( .A1(n57), .A2(pipe6_divisor_n[1]), .A3(pipe6_divisor_n[19]), 
        .ZN(n54) );
  NAND3_X1 U424 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n57) );
  NOR3_X1 U425 ( .A1(n58), .A2(pipe6_divisor_n[15]), .A3(pipe6_divisor_n[14]), 
        .ZN(n53) );
  NAND3_X1 U426 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n58) );
  NOR3_X1 U427 ( .A1(n59), .A2(pipe6_divisor_n[10]), .A3(pipe6_divisor_n[0]), 
        .ZN(n52) );
  NAND3_X1 U428 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n59) );
  INV_X1 U429 ( .A(divisor[19]), .ZN(n226) );
  INV_X1 U430 ( .A(divisor[18]), .ZN(n227) );
  INV_X1 U431 ( .A(divisor[17]), .ZN(n228) );
  INV_X1 U432 ( .A(divisor[16]), .ZN(n229) );
  INV_X1 U433 ( .A(divisor[15]), .ZN(n230) );
  INV_X1 U434 ( .A(divisor[14]), .ZN(n231) );
  INV_X1 U435 ( .A(divisor[13]), .ZN(n232) );
  INV_X1 U436 ( .A(divisor[12]), .ZN(n233) );
  INV_X1 U437 ( .A(divisor[11]), .ZN(n234) );
  INV_X1 U438 ( .A(divisor[10]), .ZN(n235) );
  INV_X1 U439 ( .A(divisor[9]), .ZN(n236) );
  INV_X1 U440 ( .A(divisor[8]), .ZN(n237) );
  INV_X1 U441 ( .A(divisor[7]), .ZN(n238) );
  INV_X1 U442 ( .A(divisor[6]), .ZN(n239) );
  INV_X1 U443 ( .A(divisor[5]), .ZN(n240) );
  INV_X1 U444 ( .A(divisor[4]), .ZN(n241) );
  INV_X1 U445 ( .A(divisor[3]), .ZN(n242) );
  INV_X1 U446 ( .A(divisor[2]), .ZN(n243) );
  INV_X1 U447 ( .A(divisor[1]), .ZN(n244) );
  INV_X1 U448 ( .A(divisor[0]), .ZN(n245) );
  NOR2_X1 U449 ( .A1(n224), .A2(n79), .ZN(N99) );
  NOR2_X1 U450 ( .A1(n224), .A2(n80), .ZN(N98) );
  NOR2_X1 U451 ( .A1(n224), .A2(n81), .ZN(N97) );
  NOR2_X1 U452 ( .A1(n224), .A2(n82), .ZN(N96) );
  NOR2_X1 U453 ( .A1(n224), .A2(n83), .ZN(N95) );
  AND2_X1 U454 ( .A1(stage1_result[27]), .A2(StartOut0), .ZN(N94) );
  AND2_X1 U455 ( .A1(stage1_result[26]), .A2(StartOut0), .ZN(N93) );
  AND2_X1 U456 ( .A1(stage1_result[25]), .A2(StartOut0), .ZN(N92) );
  AND2_X1 U457 ( .A1(stage1_result[24]), .A2(StartOut0), .ZN(N91) );
  AND2_X1 U458 ( .A1(stage1_result[23]), .A2(StartOut0), .ZN(N90) );
  AND2_X1 U459 ( .A1(stage1_result[22]), .A2(StartOut0), .ZN(N89) );
  AND2_X1 U460 ( .A1(stage1_result[21]), .A2(StartOut0), .ZN(N88) );
  AND2_X1 U461 ( .A1(stage1_result[20]), .A2(StartOut0), .ZN(N87) );
  AND2_X1 U462 ( .A1(stage1_result[19]), .A2(StartOut0), .ZN(N86) );
  AND2_X1 U463 ( .A1(stage1_result[18]), .A2(StartOut0), .ZN(N85) );
  AND2_X1 U464 ( .A1(stage1_result[17]), .A2(StartOut0), .ZN(N84) );
  AND2_X1 U465 ( .A1(stage1_result[16]), .A2(StartOut0), .ZN(N83) );
  AND2_X1 U466 ( .A1(stage1_result[15]), .A2(StartOut0), .ZN(N82) );
  AND2_X1 U467 ( .A1(stage1_result[14]), .A2(StartOut0), .ZN(N81) );
  AND2_X1 U468 ( .A1(stage1_result[13]), .A2(StartOut0), .ZN(N80) );
  AND2_X1 U469 ( .A1(stage1_result[12]), .A2(StartOut0), .ZN(N79) );
  AND2_X1 U470 ( .A1(stage1_result[11]), .A2(StartOut0), .ZN(N78) );
  AND2_X1 U471 ( .A1(stage1_result[10]), .A2(StartOut0), .ZN(N77) );
  AND2_X1 U472 ( .A1(stage1_result[9]), .A2(StartOut0), .ZN(N76) );
  AND2_X1 U473 ( .A1(stage1_result[8]), .A2(StartOut0), .ZN(N75) );
  AND2_X1 U474 ( .A1(stage1_result[7]), .A2(StartOut0), .ZN(N74) );
  AND2_X1 U475 ( .A1(stage1_result[6]), .A2(StartOut0), .ZN(N73) );
  AND2_X1 U476 ( .A1(stage1_result[5]), .A2(StartOut0), .ZN(N72) );
  AND2_X1 U477 ( .A1(stage1_result[4]), .A2(StartOut0), .ZN(N71) );
  AND2_X1 U478 ( .A1(stage1_result[3]), .A2(StartOut0), .ZN(N70) );
  AND2_X1 U479 ( .A1(stage1_result[2]), .A2(StartOut0), .ZN(N69) );
  AND2_X1 U480 ( .A1(stage1_result[1]), .A2(StartOut0), .ZN(N68) );
  AND2_X1 U481 ( .A1(start), .A2(q_bit7), .ZN(N65) );
  AND2_X1 U482 ( .A1(stage0_result[27]), .A2(start), .ZN(N44) );
  AND2_X1 U483 ( .A1(stage0_result[26]), .A2(start), .ZN(N43) );
  AND2_X1 U484 ( .A1(stage0_result[25]), .A2(start), .ZN(N42) );
  AND2_X1 U485 ( .A1(stage0_result[24]), .A2(start), .ZN(N41) );
  AND2_X1 U486 ( .A1(stage0_result[23]), .A2(start), .ZN(N40) );
  AND2_X1 U487 ( .A1(stage0_result[22]), .A2(start), .ZN(N39) );
  NOR2_X1 U488 ( .A1(n110), .A2(n84), .ZN(N386) );
  NOR2_X1 U489 ( .A1(n110), .A2(n85), .ZN(N385) );
  NOR2_X1 U490 ( .A1(n110), .A2(n86), .ZN(N384) );
  NOR2_X1 U491 ( .A1(n110), .A2(n87), .ZN(N383) );
  NOR2_X1 U492 ( .A1(n110), .A2(n88), .ZN(N382) );
  NOR2_X1 U493 ( .A1(n110), .A2(n89), .ZN(N381) );
  AND2_X1 U494 ( .A1(q_bit1), .A2(StartOut5), .ZN(N380) );
  AND2_X1 U495 ( .A1(stage0_result[21]), .A2(start), .ZN(N38) );
  NOR2_X1 U496 ( .A1(n110), .A2(n90), .ZN(N379) );
  NOR2_X1 U497 ( .A1(n110), .A2(n91), .ZN(N378) );
  NOR2_X1 U498 ( .A1(n110), .A2(n92), .ZN(N377) );
  NOR2_X1 U499 ( .A1(n110), .A2(n93), .ZN(N376) );
  NOR2_X1 U500 ( .A1(n110), .A2(n94), .ZN(N375) );
  NOR2_X1 U501 ( .A1(n110), .A2(n95), .ZN(N374) );
  NOR2_X1 U502 ( .A1(n110), .A2(n96), .ZN(N373) );
  NOR2_X1 U503 ( .A1(n110), .A2(n97), .ZN(N372) );
  NOR2_X1 U504 ( .A1(n110), .A2(n98), .ZN(N371) );
  NOR2_X1 U505 ( .A1(n110), .A2(n99), .ZN(N370) );
  AND2_X1 U506 ( .A1(stage0_result[20]), .A2(start), .ZN(N37) );
  NOR2_X1 U507 ( .A1(n110), .A2(n100), .ZN(N369) );
  NOR2_X1 U508 ( .A1(n110), .A2(n101), .ZN(N368) );
  NOR2_X1 U509 ( .A1(n110), .A2(n102), .ZN(N367) );
  NOR2_X1 U510 ( .A1(n110), .A2(n103), .ZN(N366) );
  NOR2_X1 U511 ( .A1(n110), .A2(n104), .ZN(N365) );
  NOR2_X1 U512 ( .A1(n110), .A2(n105), .ZN(N364) );
  NOR2_X1 U513 ( .A1(n110), .A2(n106), .ZN(N363) );
  NOR2_X1 U514 ( .A1(n110), .A2(n107), .ZN(N362) );
  NOR2_X1 U515 ( .A1(n110), .A2(n108), .ZN(N361) );
  NOR2_X1 U516 ( .A1(n110), .A2(n109), .ZN(N360) );
  AND2_X1 U517 ( .A1(stage0_result[19]), .A2(start), .ZN(N36) );
  AND2_X1 U518 ( .A1(stage6_result[27]), .A2(StartOut5), .ZN(N359) );
  AND2_X1 U519 ( .A1(stage6_result[26]), .A2(StartOut5), .ZN(N358) );
  AND2_X1 U520 ( .A1(stage6_result[25]), .A2(StartOut5), .ZN(N357) );
  AND2_X1 U521 ( .A1(stage6_result[24]), .A2(StartOut5), .ZN(N356) );
  AND2_X1 U522 ( .A1(stage6_result[23]), .A2(StartOut5), .ZN(N355) );
  AND2_X1 U523 ( .A1(stage6_result[22]), .A2(StartOut5), .ZN(N354) );
  AND2_X1 U524 ( .A1(stage6_result[21]), .A2(StartOut5), .ZN(N353) );
  AND2_X1 U525 ( .A1(stage6_result[20]), .A2(StartOut5), .ZN(N352) );
  AND2_X1 U526 ( .A1(stage6_result[19]), .A2(StartOut5), .ZN(N351) );
  AND2_X1 U527 ( .A1(stage6_result[18]), .A2(StartOut5), .ZN(N350) );
  AND2_X1 U528 ( .A1(stage0_result[18]), .A2(start), .ZN(N35) );
  AND2_X1 U529 ( .A1(stage6_result[17]), .A2(StartOut5), .ZN(N349) );
  AND2_X1 U530 ( .A1(stage6_result[16]), .A2(StartOut5), .ZN(N348) );
  AND2_X1 U531 ( .A1(stage6_result[15]), .A2(StartOut5), .ZN(N347) );
  AND2_X1 U532 ( .A1(stage6_result[14]), .A2(StartOut5), .ZN(N346) );
  AND2_X1 U533 ( .A1(stage6_result[13]), .A2(StartOut5), .ZN(N345) );
  AND2_X1 U534 ( .A1(stage6_result[12]), .A2(StartOut5), .ZN(N344) );
  AND2_X1 U535 ( .A1(stage6_result[11]), .A2(StartOut5), .ZN(N343) );
  AND2_X1 U536 ( .A1(stage6_result[10]), .A2(StartOut5), .ZN(N342) );
  AND2_X1 U537 ( .A1(stage6_result[9]), .A2(StartOut5), .ZN(N341) );
  AND2_X1 U538 ( .A1(stage6_result[8]), .A2(StartOut5), .ZN(N340) );
  AND2_X1 U539 ( .A1(stage0_result[17]), .A2(start), .ZN(N34) );
  AND2_X1 U540 ( .A1(stage6_result[7]), .A2(StartOut5), .ZN(N339) );
  AND2_X1 U541 ( .A1(stage6_result[6]), .A2(StartOut5), .ZN(N338) );
  AND2_X1 U542 ( .A1(stage6_result[5]), .A2(StartOut5), .ZN(N337) );
  AND2_X1 U543 ( .A1(stage6_result[4]), .A2(StartOut5), .ZN(N336) );
  AND2_X1 U544 ( .A1(stage6_result[3]), .A2(StartOut5), .ZN(N335) );
  AND2_X1 U545 ( .A1(stage6_result[2]), .A2(StartOut5), .ZN(N334) );
  AND2_X1 U546 ( .A1(stage6_result[1]), .A2(StartOut5), .ZN(N333) );
  NOR2_X1 U547 ( .A1(n136), .A2(n111), .ZN(N330) );
  AND2_X1 U548 ( .A1(stage0_result[16]), .A2(start), .ZN(N33) );
  NOR2_X1 U549 ( .A1(n136), .A2(n112), .ZN(N329) );
  NOR2_X1 U550 ( .A1(n136), .A2(n113), .ZN(N328) );
  NOR2_X1 U551 ( .A1(n136), .A2(n114), .ZN(N327) );
  NOR2_X1 U552 ( .A1(n136), .A2(n115), .ZN(N326) );
  AND2_X1 U553 ( .A1(q_bit2), .A2(StartOut4), .ZN(N325) );
  NOR2_X1 U554 ( .A1(n136), .A2(n116), .ZN(N324) );
  NOR2_X1 U555 ( .A1(n136), .A2(n117), .ZN(N323) );
  NOR2_X1 U556 ( .A1(n136), .A2(n118), .ZN(N322) );
  NOR2_X1 U557 ( .A1(n136), .A2(n119), .ZN(N321) );
  NOR2_X1 U558 ( .A1(n136), .A2(n120), .ZN(N320) );
  AND2_X1 U559 ( .A1(stage0_result[15]), .A2(start), .ZN(N32) );
  NOR2_X1 U560 ( .A1(n136), .A2(n121), .ZN(N319) );
  NOR2_X1 U561 ( .A1(n136), .A2(n122), .ZN(N318) );
  NOR2_X1 U562 ( .A1(n136), .A2(n123), .ZN(N317) );
  NOR2_X1 U563 ( .A1(n136), .A2(n124), .ZN(N316) );
  NOR2_X1 U564 ( .A1(n136), .A2(n125), .ZN(N315) );
  NOR2_X1 U565 ( .A1(n136), .A2(n126), .ZN(N314) );
  NOR2_X1 U566 ( .A1(n136), .A2(n127), .ZN(N313) );
  NOR2_X1 U567 ( .A1(n136), .A2(n128), .ZN(N312) );
  NOR2_X1 U568 ( .A1(n136), .A2(n129), .ZN(N311) );
  NOR2_X1 U569 ( .A1(n136), .A2(n130), .ZN(N310) );
  AND2_X1 U570 ( .A1(stage0_result[14]), .A2(start), .ZN(N31) );
  NOR2_X1 U571 ( .A1(n136), .A2(n131), .ZN(N309) );
  NOR2_X1 U572 ( .A1(n136), .A2(n132), .ZN(N308) );
  NOR2_X1 U573 ( .A1(n136), .A2(n133), .ZN(N307) );
  NOR2_X1 U574 ( .A1(n136), .A2(n134), .ZN(N306) );
  NOR2_X1 U575 ( .A1(n136), .A2(n135), .ZN(N305) );
  AND2_X1 U576 ( .A1(stage5_result[27]), .A2(StartOut4), .ZN(N304) );
  AND2_X1 U577 ( .A1(stage5_result[26]), .A2(StartOut4), .ZN(N303) );
  AND2_X1 U578 ( .A1(stage5_result[25]), .A2(StartOut4), .ZN(N302) );
  AND2_X1 U579 ( .A1(stage5_result[24]), .A2(StartOut4), .ZN(N301) );
  AND2_X1 U580 ( .A1(stage5_result[23]), .A2(StartOut4), .ZN(N300) );
  AND2_X1 U581 ( .A1(stage0_result[13]), .A2(start), .ZN(N30) );
  AND2_X1 U582 ( .A1(stage5_result[22]), .A2(StartOut4), .ZN(N299) );
  AND2_X1 U583 ( .A1(stage5_result[21]), .A2(StartOut4), .ZN(N298) );
  AND2_X1 U584 ( .A1(stage5_result[20]), .A2(StartOut4), .ZN(N297) );
  AND2_X1 U585 ( .A1(stage5_result[19]), .A2(StartOut4), .ZN(N296) );
  AND2_X1 U586 ( .A1(stage5_result[18]), .A2(StartOut4), .ZN(N295) );
  AND2_X1 U587 ( .A1(stage5_result[17]), .A2(StartOut4), .ZN(N294) );
  AND2_X1 U588 ( .A1(stage5_result[16]), .A2(StartOut4), .ZN(N293) );
  AND2_X1 U589 ( .A1(stage5_result[15]), .A2(StartOut4), .ZN(N292) );
  AND2_X1 U590 ( .A1(stage5_result[14]), .A2(StartOut4), .ZN(N291) );
  AND2_X1 U591 ( .A1(stage5_result[13]), .A2(StartOut4), .ZN(N290) );
  AND2_X1 U592 ( .A1(stage0_result[12]), .A2(start), .ZN(N29) );
  AND2_X1 U593 ( .A1(stage5_result[12]), .A2(StartOut4), .ZN(N289) );
  AND2_X1 U594 ( .A1(stage5_result[11]), .A2(StartOut4), .ZN(N288) );
  AND2_X1 U595 ( .A1(stage5_result[10]), .A2(StartOut4), .ZN(N287) );
  AND2_X1 U596 ( .A1(stage5_result[9]), .A2(StartOut4), .ZN(N286) );
  AND2_X1 U597 ( .A1(stage5_result[8]), .A2(StartOut4), .ZN(N285) );
  AND2_X1 U598 ( .A1(stage5_result[7]), .A2(StartOut4), .ZN(N284) );
  AND2_X1 U599 ( .A1(stage5_result[6]), .A2(StartOut4), .ZN(N283) );
  AND2_X1 U600 ( .A1(stage5_result[5]), .A2(StartOut4), .ZN(N282) );
  AND2_X1 U601 ( .A1(stage5_result[4]), .A2(StartOut4), .ZN(N281) );
  AND2_X1 U602 ( .A1(stage5_result[3]), .A2(StartOut4), .ZN(N280) );
  AND2_X1 U603 ( .A1(stage0_result[11]), .A2(start), .ZN(N28) );
  AND2_X1 U604 ( .A1(stage5_result[2]), .A2(StartOut4), .ZN(N279) );
  AND2_X1 U605 ( .A1(stage5_result[1]), .A2(StartOut4), .ZN(N278) );
  NOR2_X1 U606 ( .A1(n161), .A2(n137), .ZN(N275) );
  NOR2_X1 U607 ( .A1(n161), .A2(n138), .ZN(N274) );
  NOR2_X1 U608 ( .A1(n161), .A2(n139), .ZN(N273) );
  NOR2_X1 U609 ( .A1(n161), .A2(n140), .ZN(N272) );
  AND2_X1 U610 ( .A1(q_bit3), .A2(StartOut3), .ZN(N271) );
  NOR2_X1 U611 ( .A1(n161), .A2(n141), .ZN(N270) );
  AND2_X1 U612 ( .A1(stage0_result[10]), .A2(start), .ZN(N27) );
  NOR2_X1 U613 ( .A1(n161), .A2(n142), .ZN(N269) );
  NOR2_X1 U614 ( .A1(n161), .A2(n143), .ZN(N268) );
  NOR2_X1 U615 ( .A1(n161), .A2(n144), .ZN(N267) );
  NOR2_X1 U616 ( .A1(n161), .A2(n145), .ZN(N266) );
  NOR2_X1 U617 ( .A1(n161), .A2(n146), .ZN(N265) );
  NOR2_X1 U618 ( .A1(n161), .A2(n147), .ZN(N264) );
  NOR2_X1 U619 ( .A1(n161), .A2(n148), .ZN(N263) );
  NOR2_X1 U620 ( .A1(n161), .A2(n149), .ZN(N262) );
  NOR2_X1 U621 ( .A1(n161), .A2(n150), .ZN(N261) );
  NOR2_X1 U622 ( .A1(n161), .A2(n151), .ZN(N260) );
  AND2_X1 U623 ( .A1(stage0_result[9]), .A2(start), .ZN(N26) );
  NOR2_X1 U624 ( .A1(n161), .A2(n152), .ZN(N259) );
  NOR2_X1 U625 ( .A1(n161), .A2(n153), .ZN(N258) );
  NOR2_X1 U626 ( .A1(n161), .A2(n154), .ZN(N257) );
  NOR2_X1 U627 ( .A1(n161), .A2(n155), .ZN(N256) );
  NOR2_X1 U628 ( .A1(n161), .A2(n156), .ZN(N255) );
  NOR2_X1 U629 ( .A1(n161), .A2(n157), .ZN(N254) );
  NOR2_X1 U630 ( .A1(n161), .A2(n158), .ZN(N253) );
  NOR2_X1 U631 ( .A1(n161), .A2(n159), .ZN(N252) );
  NOR2_X1 U632 ( .A1(n161), .A2(n160), .ZN(N251) );
  AND2_X1 U633 ( .A1(stage4_result[27]), .A2(StartOut3), .ZN(N250) );
  AND2_X1 U634 ( .A1(stage0_result[8]), .A2(start), .ZN(N25) );
  AND2_X1 U635 ( .A1(stage4_result[26]), .A2(StartOut3), .ZN(N249) );
  AND2_X1 U636 ( .A1(stage4_result[25]), .A2(StartOut3), .ZN(N248) );
  AND2_X1 U637 ( .A1(stage4_result[24]), .A2(StartOut3), .ZN(N247) );
  AND2_X1 U638 ( .A1(stage4_result[23]), .A2(StartOut3), .ZN(N246) );
  AND2_X1 U639 ( .A1(stage4_result[22]), .A2(StartOut3), .ZN(N245) );
  AND2_X1 U640 ( .A1(stage4_result[21]), .A2(StartOut3), .ZN(N244) );
  AND2_X1 U641 ( .A1(stage4_result[20]), .A2(StartOut3), .ZN(N243) );
  AND2_X1 U642 ( .A1(stage4_result[19]), .A2(StartOut3), .ZN(N242) );
  AND2_X1 U643 ( .A1(stage4_result[18]), .A2(StartOut3), .ZN(N241) );
  AND2_X1 U644 ( .A1(stage4_result[17]), .A2(StartOut3), .ZN(N240) );
  AND2_X1 U645 ( .A1(stage0_result[7]), .A2(start), .ZN(N24) );
  AND2_X1 U646 ( .A1(stage4_result[16]), .A2(StartOut3), .ZN(N239) );
  AND2_X1 U647 ( .A1(stage4_result[15]), .A2(StartOut3), .ZN(N238) );
  AND2_X1 U648 ( .A1(stage4_result[14]), .A2(StartOut3), .ZN(N237) );
  AND2_X1 U649 ( .A1(stage4_result[13]), .A2(StartOut3), .ZN(N236) );
  AND2_X1 U650 ( .A1(stage4_result[12]), .A2(StartOut3), .ZN(N235) );
  AND2_X1 U651 ( .A1(stage4_result[11]), .A2(StartOut3), .ZN(N234) );
  AND2_X1 U652 ( .A1(stage4_result[10]), .A2(StartOut3), .ZN(N233) );
  AND2_X1 U653 ( .A1(stage4_result[9]), .A2(StartOut3), .ZN(N232) );
  AND2_X1 U654 ( .A1(stage4_result[8]), .A2(StartOut3), .ZN(N231) );
  AND2_X1 U655 ( .A1(stage4_result[7]), .A2(StartOut3), .ZN(N230) );
  AND2_X1 U656 ( .A1(stage0_result[6]), .A2(start), .ZN(N23) );
  AND2_X1 U657 ( .A1(stage4_result[6]), .A2(StartOut3), .ZN(N229) );
  AND2_X1 U658 ( .A1(stage4_result[5]), .A2(StartOut3), .ZN(N228) );
  AND2_X1 U659 ( .A1(stage4_result[4]), .A2(StartOut3), .ZN(N227) );
  AND2_X1 U660 ( .A1(stage4_result[3]), .A2(StartOut3), .ZN(N226) );
  AND2_X1 U661 ( .A1(stage4_result[2]), .A2(StartOut3), .ZN(N225) );
  AND2_X1 U662 ( .A1(stage4_result[1]), .A2(StartOut3), .ZN(N224) );
  NOR2_X1 U663 ( .A1(n185), .A2(n162), .ZN(N221) );
  NOR2_X1 U664 ( .A1(n185), .A2(n163), .ZN(N220) );
  AND2_X1 U665 ( .A1(stage0_result[5]), .A2(start), .ZN(N22) );
  NOR2_X1 U666 ( .A1(n185), .A2(n164), .ZN(N219) );
  AND2_X1 U667 ( .A1(q_bit4), .A2(StartOut2), .ZN(N218) );
  NOR2_X1 U668 ( .A1(n185), .A2(n165), .ZN(N217) );
  NOR2_X1 U669 ( .A1(n185), .A2(n166), .ZN(N216) );
  NOR2_X1 U670 ( .A1(n185), .A2(n167), .ZN(N215) );
  NOR2_X1 U671 ( .A1(n185), .A2(n168), .ZN(N214) );
  NOR2_X1 U672 ( .A1(n185), .A2(n169), .ZN(N213) );
  NOR2_X1 U673 ( .A1(n185), .A2(n170), .ZN(N212) );
  NOR2_X1 U674 ( .A1(n185), .A2(n171), .ZN(N211) );
  NOR2_X1 U675 ( .A1(n185), .A2(n172), .ZN(N210) );
  AND2_X1 U676 ( .A1(stage0_result[4]), .A2(start), .ZN(N21) );
  NOR2_X1 U677 ( .A1(n185), .A2(n173), .ZN(N209) );
  NOR2_X1 U678 ( .A1(n185), .A2(n174), .ZN(N208) );
  NOR2_X1 U679 ( .A1(n185), .A2(n175), .ZN(N207) );
  NOR2_X1 U680 ( .A1(n185), .A2(n176), .ZN(N206) );
  NOR2_X1 U681 ( .A1(n185), .A2(n177), .ZN(N205) );
  NOR2_X1 U682 ( .A1(n185), .A2(n178), .ZN(N204) );
  NOR2_X1 U683 ( .A1(n185), .A2(n179), .ZN(N203) );
  NOR2_X1 U684 ( .A1(n185), .A2(n180), .ZN(N202) );
  NOR2_X1 U685 ( .A1(n185), .A2(n181), .ZN(N201) );
  NOR2_X1 U686 ( .A1(n185), .A2(n182), .ZN(N200) );
  AND2_X1 U687 ( .A1(stage0_result[3]), .A2(start), .ZN(N20) );
  NOR2_X1 U688 ( .A1(n185), .A2(n183), .ZN(N199) );
  NOR2_X1 U689 ( .A1(n185), .A2(n184), .ZN(N198) );
  AND2_X1 U690 ( .A1(stage3_result[27]), .A2(StartOut2), .ZN(N197) );
  AND2_X1 U691 ( .A1(stage3_result[26]), .A2(StartOut2), .ZN(N196) );
  AND2_X1 U692 ( .A1(stage3_result[25]), .A2(StartOut2), .ZN(N195) );
  AND2_X1 U693 ( .A1(stage3_result[24]), .A2(StartOut2), .ZN(N194) );
  AND2_X1 U694 ( .A1(stage3_result[23]), .A2(StartOut2), .ZN(N193) );
  AND2_X1 U695 ( .A1(stage3_result[22]), .A2(StartOut2), .ZN(N192) );
  AND2_X1 U696 ( .A1(stage3_result[21]), .A2(StartOut2), .ZN(N191) );
  AND2_X1 U697 ( .A1(stage3_result[20]), .A2(StartOut2), .ZN(N190) );
  AND2_X1 U698 ( .A1(stage0_result[2]), .A2(start), .ZN(N19) );
  AND2_X1 U699 ( .A1(stage3_result[19]), .A2(StartOut2), .ZN(N189) );
  AND2_X1 U700 ( .A1(stage3_result[18]), .A2(StartOut2), .ZN(N188) );
  AND2_X1 U701 ( .A1(stage3_result[17]), .A2(StartOut2), .ZN(N187) );
  AND2_X1 U702 ( .A1(stage3_result[16]), .A2(StartOut2), .ZN(N186) );
  AND2_X1 U703 ( .A1(stage3_result[15]), .A2(StartOut2), .ZN(N185) );
  AND2_X1 U704 ( .A1(stage3_result[14]), .A2(StartOut2), .ZN(N184) );
  AND2_X1 U705 ( .A1(stage3_result[13]), .A2(StartOut2), .ZN(N183) );
  AND2_X1 U706 ( .A1(stage3_result[12]), .A2(StartOut2), .ZN(N182) );
  AND2_X1 U707 ( .A1(stage3_result[11]), .A2(StartOut2), .ZN(N181) );
  AND2_X1 U708 ( .A1(stage3_result[10]), .A2(StartOut2), .ZN(N180) );
  AND2_X1 U709 ( .A1(stage0_result[1]), .A2(start), .ZN(N18) );
  AND2_X1 U710 ( .A1(stage3_result[9]), .A2(StartOut2), .ZN(N179) );
  AND2_X1 U711 ( .A1(stage3_result[8]), .A2(StartOut2), .ZN(N178) );
  AND2_X1 U712 ( .A1(stage3_result[7]), .A2(StartOut2), .ZN(N177) );
  AND2_X1 U713 ( .A1(stage3_result[6]), .A2(StartOut2), .ZN(N176) );
  AND2_X1 U714 ( .A1(stage3_result[5]), .A2(StartOut2), .ZN(N175) );
  AND2_X1 U715 ( .A1(stage3_result[4]), .A2(StartOut2), .ZN(N174) );
  AND2_X1 U716 ( .A1(stage3_result[3]), .A2(StartOut2), .ZN(N173) );
  AND2_X1 U717 ( .A1(stage3_result[2]), .A2(StartOut2), .ZN(N172) );
  AND2_X1 U718 ( .A1(stage3_result[1]), .A2(StartOut2), .ZN(N171) );
  NOR2_X1 U719 ( .A1(n208), .A2(n186), .ZN(N168) );
  NOR2_X1 U720 ( .A1(n208), .A2(n187), .ZN(N167) );
  AND2_X1 U721 ( .A1(q_bit5), .A2(StartOut1), .ZN(N166) );
  NOR2_X1 U722 ( .A1(n208), .A2(n188), .ZN(N165) );
  NOR2_X1 U723 ( .A1(n208), .A2(n189), .ZN(N164) );
  NOR2_X1 U724 ( .A1(n208), .A2(n190), .ZN(N163) );
  NOR2_X1 U725 ( .A1(n208), .A2(n191), .ZN(N162) );
  NOR2_X1 U726 ( .A1(n208), .A2(n192), .ZN(N161) );
  NOR2_X1 U727 ( .A1(n208), .A2(n193), .ZN(N160) );
  NOR2_X1 U728 ( .A1(n208), .A2(n194), .ZN(N159) );
  NOR2_X1 U729 ( .A1(n208), .A2(n195), .ZN(N158) );
  NOR2_X1 U730 ( .A1(n208), .A2(n196), .ZN(N157) );
  NOR2_X1 U731 ( .A1(n208), .A2(n197), .ZN(N156) );
  NOR2_X1 U732 ( .A1(n208), .A2(n198), .ZN(N155) );
  NOR2_X1 U733 ( .A1(n208), .A2(n199), .ZN(N154) );
  NOR2_X1 U734 ( .A1(n208), .A2(n200), .ZN(N153) );
  NOR2_X1 U735 ( .A1(n208), .A2(n201), .ZN(N152) );
  NOR2_X1 U736 ( .A1(n208), .A2(n202), .ZN(N151) );
  NOR2_X1 U737 ( .A1(n208), .A2(n203), .ZN(N150) );
  NOR2_X1 U738 ( .A1(n208), .A2(n204), .ZN(N149) );
  NOR2_X1 U739 ( .A1(n208), .A2(n205), .ZN(N148) );
  NOR2_X1 U740 ( .A1(n208), .A2(n206), .ZN(N147) );
  NOR2_X1 U741 ( .A1(n208), .A2(n207), .ZN(N146) );
  AND2_X1 U742 ( .A1(stage2_result[27]), .A2(StartOut1), .ZN(N145) );
  AND2_X1 U743 ( .A1(stage2_result[26]), .A2(StartOut1), .ZN(N144) );
  AND2_X1 U744 ( .A1(stage2_result[25]), .A2(StartOut1), .ZN(N143) );
  AND2_X1 U745 ( .A1(stage2_result[24]), .A2(StartOut1), .ZN(N142) );
  AND2_X1 U746 ( .A1(stage2_result[23]), .A2(StartOut1), .ZN(N141) );
  AND2_X1 U747 ( .A1(stage2_result[22]), .A2(StartOut1), .ZN(N140) );
  AND2_X1 U748 ( .A1(stage2_result[21]), .A2(StartOut1), .ZN(N139) );
  AND2_X1 U749 ( .A1(stage2_result[20]), .A2(StartOut1), .ZN(N138) );
  AND2_X1 U750 ( .A1(stage2_result[19]), .A2(StartOut1), .ZN(N137) );
  AND2_X1 U751 ( .A1(stage2_result[18]), .A2(StartOut1), .ZN(N136) );
  AND2_X1 U752 ( .A1(stage2_result[17]), .A2(StartOut1), .ZN(N135) );
  AND2_X1 U753 ( .A1(stage2_result[16]), .A2(StartOut1), .ZN(N134) );
  AND2_X1 U754 ( .A1(stage2_result[15]), .A2(StartOut1), .ZN(N133) );
  AND2_X1 U755 ( .A1(stage2_result[14]), .A2(StartOut1), .ZN(N132) );
  AND2_X1 U756 ( .A1(stage2_result[13]), .A2(StartOut1), .ZN(N131) );
  AND2_X1 U757 ( .A1(stage2_result[12]), .A2(StartOut1), .ZN(N130) );
  AND2_X1 U758 ( .A1(stage2_result[11]), .A2(StartOut1), .ZN(N129) );
  AND2_X1 U759 ( .A1(stage2_result[10]), .A2(StartOut1), .ZN(N128) );
  AND2_X1 U760 ( .A1(stage2_result[9]), .A2(StartOut1), .ZN(N127) );
  AND2_X1 U761 ( .A1(stage2_result[8]), .A2(StartOut1), .ZN(N126) );
  AND2_X1 U762 ( .A1(stage2_result[7]), .A2(StartOut1), .ZN(N125) );
  AND2_X1 U763 ( .A1(stage2_result[6]), .A2(StartOut1), .ZN(N124) );
  AND2_X1 U764 ( .A1(stage2_result[5]), .A2(StartOut1), .ZN(N123) );
  AND2_X1 U765 ( .A1(stage2_result[4]), .A2(StartOut1), .ZN(N122) );
  AND2_X1 U766 ( .A1(stage2_result[3]), .A2(StartOut1), .ZN(N121) );
  AND2_X1 U767 ( .A1(stage2_result[2]), .A2(StartOut1), .ZN(N120) );
  AND2_X1 U768 ( .A1(stage2_result[1]), .A2(StartOut1), .ZN(N119) );
  NOR2_X1 U769 ( .A1(n224), .A2(n209), .ZN(N116) );
  AND2_X1 U770 ( .A1(q_bit6), .A2(StartOut0), .ZN(N115) );
  NOR2_X1 U771 ( .A1(n224), .A2(n210), .ZN(N114) );
  NOR2_X1 U772 ( .A1(n224), .A2(n211), .ZN(N113) );
  NOR2_X1 U773 ( .A1(n224), .A2(n212), .ZN(N112) );
  NOR2_X1 U774 ( .A1(n224), .A2(n213), .ZN(N111) );
  NOR2_X1 U775 ( .A1(n224), .A2(n214), .ZN(N110) );
  NOR2_X1 U776 ( .A1(n224), .A2(n215), .ZN(N109) );
  NOR2_X1 U777 ( .A1(n224), .A2(n216), .ZN(N108) );
  NOR2_X1 U778 ( .A1(n224), .A2(n217), .ZN(N107) );
  NOR2_X1 U779 ( .A1(n224), .A2(n218), .ZN(N106) );
  NOR2_X1 U780 ( .A1(n224), .A2(n219), .ZN(N105) );
  NOR2_X1 U781 ( .A1(n224), .A2(n220), .ZN(N104) );
  NOR2_X1 U782 ( .A1(n224), .A2(n221), .ZN(N103) );
  NOR2_X1 U783 ( .A1(n224), .A2(n222), .ZN(N102) );
  NOR2_X1 U784 ( .A1(n224), .A2(n223), .ZN(N101) );
  NOR2_X1 U785 ( .A1(n224), .A2(n225), .ZN(N100) );
endmodule



module Output_Fetch_MEM ( clock, reset_n, start, ReadBus, ReadAddress, DataOut, 
        StartOut, output_base_offset, done );
  input [127:0] ReadBus;
  output [15:0] ReadAddress;
  output [15:0] DataOut;
  input clock, reset_n, start, output_base_offset;
  output StartOut, done;
  wire   \U3/U1/DATA2_15 , \U18/Z_0 , \U18/DATA1_0 , \U17/Z_0 , \U17/DATA1_0 ,
         \U16/Z_0 , \U16/DATA1_0 , \U15/Z_0 , \U15/DATA1_0 , \U14/Z_0 ,
         \U14/DATA1_0 , \U13/Z_0 , \U13/DATA1_0 , \U12/Z_0 , \U12/DATA1_0 ,
         \U11/Z_0 , \U11/DATA1_0 , \U10/Z_0 , \U10/DATA1_0 , \U9/Z_0 ,
         \U9/DATA1_0 , \U8/Z_0 , \U8/DATA1_0 , \U7/Z_0 , \U7/DATA1_0 ,
         \U6/Z_0 , \U6/Z_1 , \U6/Z_2 , \U6/Z_3 , \U6/Z_4 , \U6/Z_5 , \U6/Z_6 ,
         \U6/Z_7 , \U6/Z_8 , \U6/Z_9 , \U6/Z_10 , \U6/Z_11 , \U6/Z_12 ,
         \U6/Z_13 , \U6/Z_14 , \U6/Z_15 , \U6/Z_16 , \U6/Z_17 , \U6/Z_18 ,
         \U6/Z_19 , \U6/Z_20 , \U6/Z_21 , \U6/Z_22 , \U6/Z_23 , \U6/Z_24 ,
         \U6/Z_25 , \U6/Z_26 , \U6/Z_27 , \U6/Z_28 , \U6/Z_29 , \U6/Z_30 ,
         \U6/Z_31 , \U6/Z_32 , \U6/Z_33 , \U6/Z_34 , \U6/Z_35 , \U6/Z_36 ,
         \U6/Z_37 , \U6/Z_38 , \U6/Z_39 , \U6/Z_40 , \U6/Z_41 , \U6/Z_42 ,
         \U6/Z_43 , \U6/Z_44 , \U6/Z_45 , \U6/Z_46 , \U6/Z_47 , \U6/Z_48 ,
         \U6/Z_49 , \U6/Z_50 , \U6/Z_51 , \U6/Z_52 , \U6/Z_53 , \U6/Z_54 ,
         \U6/Z_55 , \U6/Z_56 , \U6/Z_57 , \U6/Z_58 , \U6/Z_59 , \U6/Z_60 ,
         \U6/Z_61 , \U6/Z_62 , \U6/Z_63 , \U6/Z_64 , \U6/Z_65 , \U6/Z_66 ,
         \U6/Z_67 , \U6/Z_68 , \U6/Z_69 , \U6/Z_70 , \U6/Z_71 , \U6/Z_72 ,
         \U6/Z_73 , \U6/Z_74 , \U6/Z_75 , \U6/Z_76 , \U6/Z_77 , \U6/Z_78 ,
         \U6/Z_79 , \U6/Z_80 , \U6/Z_81 , \U6/Z_82 , \U6/Z_83 , \U6/Z_84 ,
         \U6/Z_85 , \U6/Z_86 , \U6/Z_87 , \U6/Z_88 , \U6/Z_89 , \U6/Z_90 ,
         \U6/Z_91 , \U6/Z_92 , \U6/Z_93 , \U6/Z_94 , \U6/Z_95 , \U6/Z_96 ,
         \U6/Z_97 , \U6/Z_98 , \U6/Z_99 , \U6/Z_100 , \U6/Z_101 , \U6/Z_102 ,
         \U6/Z_103 , \U6/Z_104 , \U6/Z_105 , \U6/Z_106 , \U6/Z_107 ,
         \U6/Z_108 , \U6/Z_109 , \U6/Z_110 , \U6/Z_111 , \U6/Z_112 ,
         \U6/Z_113 , \U6/Z_114 , \U6/Z_115 , \U6/Z_116 , \U6/Z_117 ,
         \U6/Z_118 , \U6/Z_119 , \U6/Z_120 , \U6/Z_121 , \U6/Z_122 ,
         \U6/Z_123 , \U6/Z_124 , \U6/Z_125 , \U6/Z_126 , \U6/Z_127 ,
         \U6/DATA2_0 , \U6/DATA2_1 , \U6/DATA2_2 , \U6/DATA2_3 , \U6/DATA2_4 ,
         \U6/DATA2_5 , \U6/DATA2_6 , \U6/DATA2_7 , \U6/DATA2_8 , \U6/DATA2_9 ,
         \U6/DATA2_10 , \U6/DATA2_11 , \U6/DATA2_12 , \U6/DATA2_13 ,
         \U6/DATA2_14 , \U6/DATA2_15 , \U6/DATA2_16 , \U6/DATA2_17 ,
         \U6/DATA2_18 , \U6/DATA2_19 , \U6/DATA2_20 , \U6/DATA2_21 ,
         \U6/DATA2_22 , \U6/DATA2_23 , \U6/DATA2_24 , \U6/DATA2_25 ,
         \U6/DATA2_26 , \U6/DATA2_27 , \U6/DATA2_28 , \U6/DATA2_29 ,
         \U6/DATA2_30 , \U6/DATA2_31 , \U6/DATA2_32 , \U6/DATA2_33 ,
         \U6/DATA2_34 , \U6/DATA2_35 , \U6/DATA2_36 , \U6/DATA2_37 ,
         \U6/DATA2_38 , \U6/DATA2_39 , \U6/DATA2_40 , \U6/DATA2_41 ,
         \U6/DATA2_42 , \U6/DATA2_43 , \U6/DATA2_44 , \U6/DATA2_45 ,
         \U6/DATA2_46 , \U6/DATA2_47 , \U6/DATA2_48 , \U6/DATA2_49 ,
         \U6/DATA2_50 , \U6/DATA2_51 , \U6/DATA2_52 , \U6/DATA2_53 ,
         \U6/DATA2_54 , \U6/DATA2_55 , \U6/DATA2_56 , \U6/DATA2_57 ,
         \U6/DATA2_58 , \U6/DATA2_59 , \U6/DATA2_60 , \U6/DATA2_61 ,
         \U6/DATA2_62 , \U6/DATA2_63 , \U6/DATA2_64 , \U6/DATA2_65 ,
         \U6/DATA2_66 , \U6/DATA2_67 , \U6/DATA2_68 , \U6/DATA2_69 ,
         \U6/DATA2_70 , \U6/DATA2_71 , \U6/DATA2_72 , \U6/DATA2_73 ,
         \U6/DATA2_74 , \U6/DATA2_75 , \U6/DATA2_76 , \U6/DATA2_77 ,
         \U6/DATA2_78 , \U6/DATA2_79 , \U6/DATA2_80 , \U6/DATA2_81 ,
         \U6/DATA2_82 , \U6/DATA2_83 , \U6/DATA2_84 , \U6/DATA2_85 ,
         \U6/DATA2_86 , \U6/DATA2_87 , \U6/DATA2_88 , \U6/DATA2_89 ,
         \U6/DATA2_90 , \U6/DATA2_91 , \U6/DATA2_92 , \U6/DATA2_93 ,
         \U6/DATA2_94 , \U6/DATA2_95 , \U6/DATA2_96 , \U6/DATA2_97 ,
         \U6/DATA2_98 , \U6/DATA2_99 , \U6/DATA2_100 , \U6/DATA2_101 ,
         \U6/DATA2_102 , \U6/DATA2_103 , \U6/DATA2_104 , \U6/DATA2_105 ,
         \U6/DATA2_106 , \U6/DATA2_107 , \U6/DATA2_108 , \U6/DATA2_109 ,
         \U6/DATA2_110 , \U6/DATA2_111 , \U6/DATA2_112 , \U6/DATA2_113 ,
         \U6/DATA2_114 , \U6/DATA2_115 , \U6/DATA2_116 , \U6/DATA2_117 ,
         \U6/DATA2_118 , \U6/DATA2_119 , \U6/DATA2_120 , \U6/DATA2_121 ,
         \U6/DATA2_122 , \U6/DATA2_123 , \U6/DATA2_124 , \U6/DATA2_125 ,
         \U6/DATA2_126 , \U6/DATA2_127 , \U5/Z_0 , \U5/Z_1 , \U5/Z_2 ,
         \U5/Z_3 , \U5/Z_4 , \U5/Z_5 , \U5/Z_6 , \U5/Z_7 , \U5/DATA16_0 ,
         \U5/DATA16_1 , \U5/DATA16_2 , \U5/DATA16_3 , \U5/DATA16_4 ,
         \U5/DATA16_5 , \U5/DATA16_6 , \U5/DATA16_7 , \U5/DATA15_0 ,
         \U5/DATA15_1 , \U5/DATA15_2 , \U5/DATA15_3 , \U5/DATA15_4 ,
         \U5/DATA15_5 , \U5/DATA15_6 , \U5/DATA15_7 , \U5/DATA14_0 ,
         \U5/DATA14_1 , \U5/DATA14_2 , \U5/DATA14_3 , \U5/DATA14_4 ,
         \U5/DATA14_5 , \U5/DATA14_6 , \U5/DATA14_7 , \U5/DATA13_0 ,
         \U5/DATA13_1 , \U5/DATA13_2 , \U5/DATA13_3 , \U5/DATA13_4 ,
         \U5/DATA13_5 , \U5/DATA13_6 , \U5/DATA13_7 , \U5/DATA12_0 ,
         \U5/DATA12_1 , \U5/DATA12_2 , \U5/DATA12_3 , \U5/DATA12_4 ,
         \U5/DATA12_5 , \U5/DATA12_6 , \U5/DATA12_7 , \U5/DATA11_0 ,
         \U5/DATA11_1 , \U5/DATA11_2 , \U5/DATA11_3 , \U5/DATA11_4 ,
         \U5/DATA11_5 , \U5/DATA11_6 , \U5/DATA11_7 , \U5/DATA10_0 ,
         \U5/DATA10_1 , \U5/DATA10_2 , \U5/DATA10_3 , \U5/DATA10_4 ,
         \U5/DATA10_5 , \U5/DATA10_6 , \U5/DATA10_7 , \U5/DATA9_0 ,
         \U5/DATA9_1 , \U5/DATA9_2 , \U5/DATA9_3 , \U5/DATA9_4 , \U5/DATA9_5 ,
         \U5/DATA9_6 , \U5/DATA9_7 , \U5/DATA8_0 , \U5/DATA8_1 , \U5/DATA8_2 ,
         \U5/DATA8_3 , \U5/DATA8_4 , \U5/DATA8_5 , \U5/DATA8_6 , \U5/DATA8_7 ,
         \U5/DATA7_0 , \U5/DATA7_1 , \U5/DATA7_2 , \U5/DATA7_3 , \U5/DATA7_4 ,
         \U5/DATA7_5 , \U5/DATA7_6 , \U5/DATA7_7 , \U5/DATA6_0 , \U5/DATA6_1 ,
         \U5/DATA6_2 , \U5/DATA6_3 , \U5/DATA6_4 , \U5/DATA6_5 , \U5/DATA6_6 ,
         \U5/DATA6_7 , \U5/DATA5_0 , \U5/DATA5_1 , \U5/DATA5_2 , \U5/DATA5_3 ,
         \U5/DATA5_4 , \U5/DATA5_5 , \U5/DATA5_6 , \U5/DATA5_7 , \U5/DATA4_0 ,
         \U5/DATA4_1 , \U5/DATA4_2 , \U5/DATA4_3 , \U5/DATA4_4 , \U5/DATA4_5 ,
         \U5/DATA4_6 , \U5/DATA4_7 , \U5/DATA3_0 , \U5/DATA3_1 , \U5/DATA3_2 ,
         \U5/DATA3_3 , \U5/DATA3_4 , \U5/DATA3_5 , \U5/DATA3_6 , \U5/DATA3_7 ,
         \U5/DATA2_0 , \U5/DATA2_1 , \U5/DATA2_2 , \U5/DATA2_3 , \U5/DATA2_4 ,
         \U5/DATA2_5 , \U5/DATA2_6 , \U5/DATA2_7 , \U5/DATA1_0 , \U5/DATA1_1 ,
         \U5/DATA1_2 , \U5/DATA1_3 , \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 ,
         \U5/DATA1_7 , \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \add_101/A[0] ,
         \add_101/A[1] , \add_101/A[2] , \add_101/A[3] , \add_101/A[4] ,
         \add_101/A[5] , \add_101/A[6] , \add_101/A[7] , \add_101/A[8] ,
         \add_101/A[9] , \add_101/A[10] , \add_101/A[11] , \add_101/A[12] ,
         \add_101/A[13] , \add_101/A[14] , \add_101/A[15] , \add_95/A[0] ,
         \add_95/A[1] , \add_95/A[2] , \add_95/A[3] , n22, n24, n25, n26, n27,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n147, n148,
         n149, n150, n151, n153, n154, n155, n156, n161, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739;
  assign \U3/U1/DATA2_15  = output_base_offset;
  assign \U6/DATA2_0  = ReadBus[0];
  assign \U6/DATA2_1  = ReadBus[1];
  assign \U6/DATA2_2  = ReadBus[2];
  assign \U6/DATA2_3  = ReadBus[3];
  assign \U6/DATA2_4  = ReadBus[4];
  assign \U6/DATA2_5  = ReadBus[5];
  assign \U6/DATA2_6  = ReadBus[6];
  assign \U6/DATA2_7  = ReadBus[7];
  assign \U6/DATA2_8  = ReadBus[8];
  assign \U6/DATA2_9  = ReadBus[9];
  assign \U6/DATA2_10  = ReadBus[10];
  assign \U6/DATA2_11  = ReadBus[11];
  assign \U6/DATA2_12  = ReadBus[12];
  assign \U6/DATA2_13  = ReadBus[13];
  assign \U6/DATA2_14  = ReadBus[14];
  assign \U6/DATA2_15  = ReadBus[15];
  assign \U6/DATA2_16  = ReadBus[16];
  assign \U6/DATA2_17  = ReadBus[17];
  assign \U6/DATA2_18  = ReadBus[18];
  assign \U6/DATA2_19  = ReadBus[19];
  assign \U6/DATA2_20  = ReadBus[20];
  assign \U6/DATA2_21  = ReadBus[21];
  assign \U6/DATA2_22  = ReadBus[22];
  assign \U6/DATA2_23  = ReadBus[23];
  assign \U6/DATA2_24  = ReadBus[24];
  assign \U6/DATA2_25  = ReadBus[25];
  assign \U6/DATA2_26  = ReadBus[26];
  assign \U6/DATA2_27  = ReadBus[27];
  assign \U6/DATA2_28  = ReadBus[28];
  assign \U6/DATA2_29  = ReadBus[29];
  assign \U6/DATA2_30  = ReadBus[30];
  assign \U6/DATA2_31  = ReadBus[31];
  assign \U6/DATA2_32  = ReadBus[32];
  assign \U6/DATA2_33  = ReadBus[33];
  assign \U6/DATA2_34  = ReadBus[34];
  assign \U6/DATA2_35  = ReadBus[35];
  assign \U6/DATA2_36  = ReadBus[36];
  assign \U6/DATA2_37  = ReadBus[37];
  assign \U6/DATA2_38  = ReadBus[38];
  assign \U6/DATA2_39  = ReadBus[39];
  assign \U6/DATA2_40  = ReadBus[40];
  assign \U6/DATA2_41  = ReadBus[41];
  assign \U6/DATA2_42  = ReadBus[42];
  assign \U6/DATA2_43  = ReadBus[43];
  assign \U6/DATA2_44  = ReadBus[44];
  assign \U6/DATA2_45  = ReadBus[45];
  assign \U6/DATA2_46  = ReadBus[46];
  assign \U6/DATA2_47  = ReadBus[47];
  assign \U6/DATA2_48  = ReadBus[48];
  assign \U6/DATA2_49  = ReadBus[49];
  assign \U6/DATA2_50  = ReadBus[50];
  assign \U6/DATA2_51  = ReadBus[51];
  assign \U6/DATA2_52  = ReadBus[52];
  assign \U6/DATA2_53  = ReadBus[53];
  assign \U6/DATA2_54  = ReadBus[54];
  assign \U6/DATA2_55  = ReadBus[55];
  assign \U6/DATA2_56  = ReadBus[56];
  assign \U6/DATA2_57  = ReadBus[57];
  assign \U6/DATA2_58  = ReadBus[58];
  assign \U6/DATA2_59  = ReadBus[59];
  assign \U6/DATA2_60  = ReadBus[60];
  assign \U6/DATA2_61  = ReadBus[61];
  assign \U6/DATA2_62  = ReadBus[62];
  assign \U6/DATA2_63  = ReadBus[63];
  assign \U6/DATA2_64  = ReadBus[64];
  assign \U6/DATA2_65  = ReadBus[65];
  assign \U6/DATA2_66  = ReadBus[66];
  assign \U6/DATA2_67  = ReadBus[67];
  assign \U6/DATA2_68  = ReadBus[68];
  assign \U6/DATA2_69  = ReadBus[69];
  assign \U6/DATA2_70  = ReadBus[70];
  assign \U6/DATA2_71  = ReadBus[71];
  assign \U6/DATA2_72  = ReadBus[72];
  assign \U6/DATA2_73  = ReadBus[73];
  assign \U6/DATA2_74  = ReadBus[74];
  assign \U6/DATA2_75  = ReadBus[75];
  assign \U6/DATA2_76  = ReadBus[76];
  assign \U6/DATA2_77  = ReadBus[77];
  assign \U6/DATA2_78  = ReadBus[78];
  assign \U6/DATA2_79  = ReadBus[79];
  assign \U6/DATA2_80  = ReadBus[80];
  assign \U6/DATA2_81  = ReadBus[81];
  assign \U6/DATA2_82  = ReadBus[82];
  assign \U6/DATA2_83  = ReadBus[83];
  assign \U6/DATA2_84  = ReadBus[84];
  assign \U6/DATA2_85  = ReadBus[85];
  assign \U6/DATA2_86  = ReadBus[86];
  assign \U6/DATA2_87  = ReadBus[87];
  assign \U6/DATA2_88  = ReadBus[88];
  assign \U6/DATA2_89  = ReadBus[89];
  assign \U6/DATA2_90  = ReadBus[90];
  assign \U6/DATA2_91  = ReadBus[91];
  assign \U6/DATA2_92  = ReadBus[92];
  assign \U6/DATA2_93  = ReadBus[93];
  assign \U6/DATA2_94  = ReadBus[94];
  assign \U6/DATA2_95  = ReadBus[95];
  assign \U6/DATA2_96  = ReadBus[96];
  assign \U6/DATA2_97  = ReadBus[97];
  assign \U6/DATA2_98  = ReadBus[98];
  assign \U6/DATA2_99  = ReadBus[99];
  assign \U6/DATA2_100  = ReadBus[100];
  assign \U6/DATA2_101  = ReadBus[101];
  assign \U6/DATA2_102  = ReadBus[102];
  assign \U6/DATA2_103  = ReadBus[103];
  assign \U6/DATA2_104  = ReadBus[104];
  assign \U6/DATA2_105  = ReadBus[105];
  assign \U6/DATA2_106  = ReadBus[106];
  assign \U6/DATA2_107  = ReadBus[107];
  assign \U6/DATA2_108  = ReadBus[108];
  assign \U6/DATA2_109  = ReadBus[109];
  assign \U6/DATA2_110  = ReadBus[110];
  assign \U6/DATA2_111  = ReadBus[111];
  assign \U6/DATA2_112  = ReadBus[112];
  assign \U6/DATA2_113  = ReadBus[113];
  assign \U6/DATA2_114  = ReadBus[114];
  assign \U6/DATA2_115  = ReadBus[115];
  assign \U6/DATA2_116  = ReadBus[116];
  assign \U6/DATA2_117  = ReadBus[117];
  assign \U6/DATA2_118  = ReadBus[118];
  assign \U6/DATA2_119  = ReadBus[119];
  assign \U6/DATA2_120  = ReadBus[120];
  assign \U6/DATA2_121  = ReadBus[121];
  assign \U6/DATA2_122  = ReadBus[122];
  assign \U6/DATA2_123  = ReadBus[123];
  assign \U6/DATA2_124  = ReadBus[124];
  assign \U6/DATA2_125  = ReadBus[125];
  assign \U6/DATA2_126  = ReadBus[126];
  assign \U6/DATA2_127  = ReadBus[127];
  assign DataOut[0] = \U5/Z_0 ;
  assign DataOut[1] = \U5/Z_1 ;
  assign DataOut[2] = \U5/Z_2 ;
  assign DataOut[3] = \U5/Z_3 ;
  assign DataOut[4] = \U5/Z_4 ;
  assign DataOut[5] = \U5/Z_5 ;
  assign DataOut[6] = \U5/Z_6 ;
  assign DataOut[7] = \U5/Z_7 ;
  assign ReadAddress[0] = \add_101/A[0] ;
  assign ReadAddress[1] = \add_101/A[1] ;
  assign ReadAddress[2] = \add_101/A[2] ;
  assign ReadAddress[3] = \add_101/A[3] ;
  assign ReadAddress[4] = \add_101/A[4] ;
  assign ReadAddress[5] = \add_101/A[5] ;
  assign ReadAddress[6] = \add_101/A[6] ;
  assign ReadAddress[7] = \add_101/A[7] ;
  assign ReadAddress[8] = \add_101/A[8] ;
  assign ReadAddress[9] = \add_101/A[9] ;
  assign ReadAddress[10] = \add_101/A[10] ;
  assign ReadAddress[11] = \add_101/A[11] ;
  assign ReadAddress[12] = \add_101/A[12] ;
  assign ReadAddress[13] = \add_101/A[13] ;
  assign ReadAddress[14] = \add_101/A[14] ;
  assign ReadAddress[15] = \add_101/A[15] ;

  DFFR_X1 \short_count_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n632), .Q(
        \add_95/A[0] ), .QN(n27) );
  DFFR_X1 \short_count_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .RN(n628), .Q(
        \add_95/A[2] ), .QN(n25) );
  DFFR_X1 \short_count_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n628), .Q(
        \add_95/A[3] ), .QN(n24) );
  DFFR_X1 done0_reg ( .D(n739), .CK(clock), .RN(n629), .Q(\U18/DATA1_0 ) );
  DFFR_X1 done1_reg ( .D(\U18/Z_0 ), .CK(clock), .RN(n629), .Q(\U17/DATA1_0 )
         );
  DFFR_X1 done2_reg ( .D(\U17/Z_0 ), .CK(clock), .RN(n629), .Q(\U16/DATA1_0 )
         );
  DFFR_X1 done3_reg ( .D(\U16/Z_0 ), .CK(clock), .RN(n629), .Q(\U15/DATA1_0 )
         );
  DFFR_X1 done4_reg ( .D(\U15/Z_0 ), .CK(clock), .RN(n629), .Q(\U14/DATA1_0 )
         );
  DFFR_X1 done5_reg ( .D(\U14/Z_0 ), .CK(clock), .RN(n636), .Q(\U13/DATA1_0 )
         );
  DFFR_X1 done6_reg ( .D(\U13/Z_0 ), .CK(clock), .RN(n637), .Q(\U12/DATA1_0 )
         );
  DFFR_X1 done7_reg ( .D(\U12/Z_0 ), .CK(clock), .RN(n637), .Q(\U11/DATA1_0 )
         );
  DFFR_X1 done8_reg ( .D(\U11/Z_0 ), .CK(clock), .RN(n637), .Q(\U10/DATA1_0 )
         );
  DFFR_X1 done9_reg ( .D(\U10/Z_0 ), .CK(clock), .RN(n637), .Q(\U9/DATA1_0 )
         );
  DFFR_X1 done10_reg ( .D(\U9/Z_0 ), .CK(clock), .RN(n637), .Q(\U8/DATA1_0 )
         );
  DFFR_X1 done11_reg ( .D(\U8/Z_0 ), .CK(clock), .RN(n637), .Q(\U7/DATA1_0 )
         );
  DFFR_X1 done_reg ( .D(\U7/Z_0 ), .CK(clock), .RN(n637), .Q(done) );
  SDFFR_X2 StartOut_reg ( .D(1'b0), .SI(n50), .SE(start), .CK(clock), .RN(n637), .Q(StartOut) );
  DFFR_X1 \data_in_reg[0]  ( .D(\U6/Z_0 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA16_0 ) );
  DFFR_X1 \data_in_reg[1]  ( .D(\U6/Z_1 ), .CK(clock), .RN(n637), .Q(
        \U5/DATA16_1 ) );
  DFFR_X1 \data_in_reg[10]  ( .D(\U6/Z_10 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA1_2 ) );
  DFFR_X1 \data_in_reg[100]  ( .D(\U6/Z_100 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA12_4 ) );
  DFFR_X1 \data_in_reg[101]  ( .D(\U6/Z_101 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA12_5 ) );
  DFFR_X1 \data_in_reg[102]  ( .D(\U6/Z_102 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA12_6 ) );
  DFFR_X1 \data_in_reg[103]  ( .D(\U6/Z_103 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA12_7 ) );
  DFFR_X1 \data_in_reg[104]  ( .D(\U6/Z_104 ), .CK(clock), .RN(n637), .Q(
        \U5/DATA13_0 ) );
  DFFR_X1 \data_in_reg[105]  ( .D(\U6/Z_105 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA13_1 ) );
  DFFR_X1 \data_in_reg[106]  ( .D(\U6/Z_106 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA13_2 ) );
  DFFR_X1 \data_in_reg[107]  ( .D(\U6/Z_107 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA13_3 ) );
  DFFR_X1 \data_in_reg[108]  ( .D(\U6/Z_108 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA13_4 ) );
  DFFR_X1 \data_in_reg[109]  ( .D(\U6/Z_109 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA13_5 ) );
  DFFR_X1 \data_in_reg[11]  ( .D(\U6/Z_11 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA1_3 ) );
  DFFR_X1 \data_in_reg[110]  ( .D(\U6/Z_110 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA13_6 ) );
  DFFR_X1 \data_in_reg[111]  ( .D(\U6/Z_111 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA13_7 ) );
  DFFR_X1 \data_in_reg[112]  ( .D(\U6/Z_112 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA14_0 ) );
  DFFR_X1 \data_in_reg[113]  ( .D(\U6/Z_113 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA14_1 ) );
  DFFR_X1 \data_in_reg[114]  ( .D(\U6/Z_114 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA14_2 ) );
  DFFR_X1 \data_in_reg[115]  ( .D(\U6/Z_115 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA14_3 ) );
  DFFR_X1 \data_in_reg[116]  ( .D(\U6/Z_116 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA14_4 ) );
  DFFR_X1 \data_in_reg[117]  ( .D(\U6/Z_117 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA14_5 ) );
  DFFR_X1 \data_in_reg[118]  ( .D(\U6/Z_118 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA14_6 ) );
  DFFR_X1 \data_in_reg[119]  ( .D(\U6/Z_119 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA14_7 ) );
  DFFR_X1 \data_in_reg[12]  ( .D(\U6/Z_12 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA1_4 ) );
  DFFR_X1 \data_in_reg[120]  ( .D(\U6/Z_120 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA15_0 ) );
  DFFR_X1 \data_in_reg[121]  ( .D(\U6/Z_121 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA15_1 ) );
  DFFR_X1 \data_in_reg[122]  ( .D(\U6/Z_122 ), .CK(clock), .RN(n630), .Q(
        \U5/DATA15_2 ) );
  DFFR_X1 \data_in_reg[123]  ( .D(\U6/Z_123 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA15_3 ) );
  DFFR_X1 \data_in_reg[124]  ( .D(\U6/Z_124 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA15_4 ) );
  DFFR_X1 \data_in_reg[125]  ( .D(\U6/Z_125 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA15_5 ) );
  DFFR_X1 \data_in_reg[126]  ( .D(\U6/Z_126 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA15_6 ) );
  DFFR_X1 \data_in_reg[127]  ( .D(\U6/Z_127 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA15_7 ) );
  DFFR_X1 \data_in_reg[13]  ( .D(\U6/Z_13 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA1_5 ) );
  DFFR_X1 \data_in_reg[14]  ( .D(\U6/Z_14 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA1_6 ) );
  DFFR_X1 \data_in_reg[15]  ( .D(\U6/Z_15 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA1_7 ) );
  DFFR_X1 \data_in_reg[16]  ( .D(\U6/Z_16 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA2_0 ) );
  DFFR_X1 \data_in_reg[17]  ( .D(\U6/Z_17 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA2_1 ) );
  DFFR_X1 \data_in_reg[18]  ( .D(\U6/Z_18 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA2_2 ) );
  DFFR_X1 \data_in_reg[19]  ( .D(\U6/Z_19 ), .CK(clock), .RN(n631), .Q(
        \U5/DATA2_3 ) );
  DFFR_X1 \data_in_reg[2]  ( .D(\U6/Z_2 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA16_2 ) );
  DFFR_X1 \data_in_reg[20]  ( .D(\U6/Z_20 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA2_4 ) );
  DFFR_X1 \data_in_reg[21]  ( .D(\U6/Z_21 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA2_5 ) );
  DFFR_X1 \data_in_reg[22]  ( .D(\U6/Z_22 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA2_6 ) );
  DFFR_X1 \data_in_reg[23]  ( .D(\U6/Z_23 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA2_7 ) );
  DFFR_X1 \data_in_reg[24]  ( .D(\U6/Z_24 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA3_0 ) );
  DFFR_X1 \data_in_reg[25]  ( .D(\U6/Z_25 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA3_1 ) );
  DFFR_X1 \data_in_reg[26]  ( .D(\U6/Z_26 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA3_2 ) );
  DFFR_X1 \data_in_reg[27]  ( .D(\U6/Z_27 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA3_3 ) );
  DFFR_X1 \data_in_reg[28]  ( .D(\U6/Z_28 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA3_4 ) );
  DFFR_X1 \data_in_reg[29]  ( .D(\U6/Z_29 ), .CK(clock), .RN(n632), .Q(
        \U5/DATA3_5 ) );
  DFFR_X1 \data_in_reg[3]  ( .D(\U6/Z_3 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA16_3 ) );
  DFFR_X1 \data_in_reg[30]  ( .D(\U6/Z_30 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA3_6 ) );
  DFFR_X1 \data_in_reg[31]  ( .D(\U6/Z_31 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA3_7 ) );
  DFFR_X1 \data_in_reg[32]  ( .D(\U6/Z_32 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA4_0 ) );
  DFFR_X1 \data_in_reg[33]  ( .D(\U6/Z_33 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA4_1 ) );
  DFFR_X1 \data_in_reg[34]  ( .D(\U6/Z_34 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA4_2 ) );
  DFFR_X1 \data_in_reg[35]  ( .D(\U6/Z_35 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA4_3 ) );
  DFFR_X1 \data_in_reg[36]  ( .D(\U6/Z_36 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA4_4 ) );
  DFFR_X1 \data_in_reg[37]  ( .D(\U6/Z_37 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA4_5 ) );
  DFFR_X1 \data_in_reg[38]  ( .D(\U6/Z_38 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA4_6 ) );
  DFFR_X1 \data_in_reg[39]  ( .D(\U6/Z_39 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA4_7 ) );
  DFFR_X1 \data_in_reg[4]  ( .D(\U6/Z_4 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA16_4 ) );
  DFFR_X1 \data_in_reg[40]  ( .D(\U6/Z_40 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA5_0 ) );
  DFFR_X1 \data_in_reg[41]  ( .D(\U6/Z_41 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA5_1 ) );
  DFFR_X1 \data_in_reg[42]  ( .D(\U6/Z_42 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA5_2 ) );
  DFFR_X1 \data_in_reg[43]  ( .D(\U6/Z_43 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA5_3 ) );
  DFFR_X1 \data_in_reg[44]  ( .D(\U6/Z_44 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA5_4 ) );
  DFFR_X1 \data_in_reg[45]  ( .D(\U6/Z_45 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA5_5 ) );
  DFFR_X1 \data_in_reg[46]  ( .D(\U6/Z_46 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA5_6 ) );
  DFFR_X1 \data_in_reg[47]  ( .D(\U6/Z_47 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA5_7 ) );
  DFFR_X1 \data_in_reg[48]  ( .D(\U6/Z_48 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA6_0 ) );
  DFFR_X1 \data_in_reg[49]  ( .D(\U6/Z_49 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA6_1 ) );
  DFFR_X1 \data_in_reg[5]  ( .D(\U6/Z_5 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA16_5 ) );
  DFFR_X1 \data_in_reg[50]  ( .D(\U6/Z_50 ), .CK(clock), .RN(n633), .Q(
        \U5/DATA6_2 ) );
  DFFR_X1 \data_in_reg[51]  ( .D(\U6/Z_51 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA6_3 ) );
  DFFR_X1 \data_in_reg[52]  ( .D(\U6/Z_52 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA6_4 ) );
  DFFR_X1 \data_in_reg[53]  ( .D(\U6/Z_53 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA6_5 ) );
  DFFR_X1 \data_in_reg[54]  ( .D(\U6/Z_54 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA6_6 ) );
  DFFR_X1 \data_in_reg[55]  ( .D(\U6/Z_55 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA6_7 ) );
  DFFR_X1 \data_in_reg[56]  ( .D(\U6/Z_56 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA7_0 ) );
  DFFR_X1 \data_in_reg[57]  ( .D(\U6/Z_57 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA7_1 ) );
  DFFR_X1 \data_in_reg[58]  ( .D(\U6/Z_58 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA7_2 ) );
  DFFR_X1 \data_in_reg[59]  ( .D(\U6/Z_59 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA7_3 ) );
  DFFR_X1 \data_in_reg[6]  ( .D(\U6/Z_6 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA16_6 ) );
  DFFR_X1 \data_in_reg[60]  ( .D(\U6/Z_60 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA7_4 ) );
  DFFR_X1 \data_in_reg[61]  ( .D(\U6/Z_61 ), .CK(clock), .RN(n634), .Q(
        \U5/DATA7_5 ) );
  DFFR_X1 \data_in_reg[62]  ( .D(\U6/Z_62 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA7_6 ) );
  DFFR_X1 \data_in_reg[63]  ( .D(\U6/Z_63 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA7_7 ) );
  DFFR_X1 \data_in_reg[64]  ( .D(\U6/Z_64 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA8_0 ) );
  DFFR_X1 \data_in_reg[65]  ( .D(\U6/Z_65 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA8_1 ) );
  DFFR_X1 \data_in_reg[66]  ( .D(\U6/Z_66 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA8_2 ) );
  DFFR_X1 \data_in_reg[67]  ( .D(\U6/Z_67 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA8_3 ) );
  DFFR_X1 \data_in_reg[68]  ( .D(\U6/Z_68 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA8_4 ) );
  DFFR_X1 \data_in_reg[69]  ( .D(\U6/Z_69 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA8_5 ) );
  DFFR_X1 \data_in_reg[7]  ( .D(\U6/Z_7 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA16_7 ) );
  DFFR_X1 \data_in_reg[70]  ( .D(\U6/Z_70 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA8_6 ) );
  DFFR_X1 \data_in_reg[71]  ( .D(\U6/Z_71 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA8_7 ) );
  DFFR_X1 \data_in_reg[72]  ( .D(\U6/Z_72 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA9_0 ) );
  DFFR_X1 \data_in_reg[73]  ( .D(\U6/Z_73 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA9_1 ) );
  DFFR_X1 \data_in_reg[74]  ( .D(\U6/Z_74 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA9_2 ) );
  DFFR_X1 \data_in_reg[75]  ( .D(\U6/Z_75 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA9_3 ) );
  DFFR_X1 \data_in_reg[76]  ( .D(\U6/Z_76 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA9_4 ) );
  DFFR_X1 \data_in_reg[77]  ( .D(\U6/Z_77 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA9_5 ) );
  DFFR_X1 \data_in_reg[78]  ( .D(\U6/Z_78 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA9_6 ) );
  DFFR_X1 \data_in_reg[79]  ( .D(\U6/Z_79 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA9_7 ) );
  DFFR_X1 \data_in_reg[8]  ( .D(\U6/Z_8 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA1_0 ) );
  DFFR_X1 \data_in_reg[80]  ( .D(\U6/Z_80 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA10_0 ) );
  DFFR_X1 \data_in_reg[81]  ( .D(\U6/Z_81 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA10_1 ) );
  DFFR_X1 \data_in_reg[82]  ( .D(\U6/Z_82 ), .CK(clock), .RN(n636), .Q(
        \U5/DATA10_2 ) );
  DFFR_X1 \data_in_reg[83]  ( .D(\U6/Z_83 ), .CK(clock), .RN(n628), .Q(
        \U5/DATA10_3 ) );
  DFFR_X1 \data_in_reg[84]  ( .D(\U6/Z_84 ), .CK(clock), .RN(n635), .Q(
        \U5/DATA10_4 ) );
  DFFR_X1 \data_in_reg[85]  ( .D(\U6/Z_85 ), .CK(clock), .RN(n629), .Q(
        \U5/DATA10_5 ) );
  DFFR_X1 \data_in_reg[86]  ( .D(\U6/Z_86 ), .CK(clock), .RN(n638), .Q(
        \U5/DATA10_6 ) );
  DFFR_X1 \data_in_reg[87]  ( .D(\U6/Z_87 ), .CK(clock), .RN(reset_n), .Q(
        \U5/DATA10_7 ) );
  DFFR_X1 \data_in_reg[88]  ( .D(\U6/Z_88 ), .CK(clock), .RN(reset_n), .Q(
        \U5/DATA11_0 ) );
  DFFR_X1 \data_in_reg[89]  ( .D(\U6/Z_89 ), .CK(clock), .RN(reset_n), .Q(
        \U5/DATA11_1 ) );
  DFFR_X1 \data_in_reg[9]  ( .D(\U6/Z_9 ), .CK(clock), .RN(reset_n), .Q(
        \U5/DATA1_1 ) );
  DFFR_X1 \data_in_reg[90]  ( .D(\U6/Z_90 ), .CK(clock), .RN(reset_n), .Q(
        \U5/DATA11_2 ) );
  DFFR_X1 \data_in_reg[91]  ( .D(\U6/Z_91 ), .CK(clock), .RN(reset_n), .Q(
        \U5/DATA11_3 ) );
  DFFR_X1 \data_in_reg[92]  ( .D(\U6/Z_92 ), .CK(clock), .RN(reset_n), .Q(
        \U5/DATA11_4 ) );
  DFFR_X1 \data_in_reg[93]  ( .D(\U6/Z_93 ), .CK(clock), .RN(n628), .Q(
        \U5/DATA11_5 ) );
  DFFR_X1 \data_in_reg[94]  ( .D(\U6/Z_94 ), .CK(clock), .RN(n637), .Q(
        \U5/DATA11_6 ) );
  DFFR_X1 \data_in_reg[95]  ( .D(\U6/Z_95 ), .CK(clock), .RN(n637), .Q(
        \U5/DATA11_7 ) );
  DFFR_X1 \data_in_reg[96]  ( .D(\U6/Z_96 ), .CK(clock), .RN(n637), .Q(
        \U5/DATA12_0 ) );
  DFFR_X1 \data_in_reg[97]  ( .D(\U6/Z_97 ), .CK(clock), .RN(n637), .Q(
        \U5/DATA12_1 ) );
  DFFR_X1 \data_in_reg[98]  ( .D(\U6/Z_98 ), .CK(clock), .RN(n637), .Q(
        \U5/DATA12_2 ) );
  DFFR_X1 \data_in_reg[99]  ( .D(\U6/Z_99 ), .CK(clock), .RN(n629), .Q(
        \U5/DATA12_3 ) );
  DFFR_X1 \short_count_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .RN(n628), .Q(
        \add_95/A[1] ), .QN(n26) );
  NAND4_X2 U25 ( .A1(n53), .A2(n54), .A3(n55), .A4(n56), .ZN(n52) );
  NAND4_X2 U30 ( .A1(n65), .A2(n66), .A3(n67), .A4(n68), .ZN(n51) );
  NAND4_X2 U35 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(n77) );
  NAND4_X2 U40 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(n76) );
  NAND4_X2 U45 ( .A1(n88), .A2(n89), .A3(n90), .A4(n91), .ZN(n87) );
  NAND4_X2 U50 ( .A1(n92), .A2(n93), .A3(n94), .A4(n95), .ZN(n86) );
  NAND4_X2 U55 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(n97) );
  NAND4_X2 U60 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(n96) );
  NAND4_X2 U65 ( .A1(n108), .A2(n109), .A3(n110), .A4(n111), .ZN(n107) );
  NAND4_X2 U70 ( .A1(n112), .A2(n113), .A3(n114), .A4(n115), .ZN(n106) );
  NAND4_X2 U75 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(n117) );
  NAND4_X2 U80 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(n116) );
  NAND4_X2 U85 ( .A1(n128), .A2(n129), .A3(n130), .A4(n131), .ZN(n127) );
  NAND4_X2 U90 ( .A1(n132), .A2(n133), .A3(n134), .A4(n135), .ZN(n126) );
  NAND4_X2 U95 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(n137) );
  NOR2_X2 U100 ( .A1(n24), .A2(\add_95/A[0] ), .ZN(n144) );
  NAND4_X2 U101 ( .A1(n148), .A2(n149), .A3(n150), .A4(n151), .ZN(n136) );
  NOR2_X2 U103 ( .A1(\add_95/A[2] ), .A2(\add_95/A[1] ), .ZN(n142) );
  NOR2_X2 U107 ( .A1(\add_95/A[3] ), .A2(\add_95/A[0] ), .ZN(n153) );
  OAI22_X2 U108 ( .A1(n154), .A2(n48), .B1(n48), .B2(n24), .ZN(\U4/Z_3 ) );
  NAND2_X2 U109 ( .A1(n625), .A2(n147), .ZN(n154) );
  OAI22_X2 U111 ( .A1(n25), .A2(n721), .B1(n155), .B2(n48), .ZN(\U4/Z_2 ) );
  NOR2_X2 U115 ( .A1(n156), .A2(n48), .ZN(\U4/Z_1 ) );
  XOR2_X2 U116 ( .A(n26), .B(\add_95/A[0] ), .Z(n156) );
  NOR2_X2 U117 ( .A1(n48), .A2(\add_95/A[0] ), .ZN(\U4/Z_0 ) );
  NAND2_X2 U118 ( .A1(n49), .A2(n50), .ZN(n48) );
  NOR2_X2 U125 ( .A1(n24), .A2(n27), .ZN(n143) );
  NOR2_X2 U126 ( .A1(n25), .A2(n26), .ZN(n147) );
  AND2_X1 U149 ( .A1(\U9/DATA1_0 ), .A2(start), .ZN(\U9/Z_0 ) );
  AND2_X1 U150 ( .A1(\U8/DATA1_0 ), .A2(start), .ZN(\U8/Z_0 ) );
  AND2_X1 U151 ( .A1(\U7/DATA1_0 ), .A2(start), .ZN(\U7/Z_0 ) );
  AND2_X1 U152 ( .A1(\U6/DATA2_99 ), .A2(n627), .ZN(\U6/Z_99 ) );
  AND2_X1 U153 ( .A1(\U6/DATA2_98 ), .A2(n626), .ZN(\U6/Z_98 ) );
  AND2_X1 U154 ( .A1(\U6/DATA2_97 ), .A2(n627), .ZN(\U6/Z_97 ) );
  AND2_X1 U155 ( .A1(\U6/DATA2_96 ), .A2(n626), .ZN(\U6/Z_96 ) );
  AND2_X1 U156 ( .A1(\U6/DATA2_95 ), .A2(n627), .ZN(\U6/Z_95 ) );
  AND2_X1 U157 ( .A1(\U6/DATA2_94 ), .A2(n627), .ZN(\U6/Z_94 ) );
  AND2_X1 U158 ( .A1(\U6/DATA2_93 ), .A2(n627), .ZN(\U6/Z_93 ) );
  AND2_X1 U159 ( .A1(\U6/DATA2_92 ), .A2(n627), .ZN(\U6/Z_92 ) );
  AND2_X1 U160 ( .A1(\U6/DATA2_91 ), .A2(n626), .ZN(\U6/Z_91 ) );
  AND2_X1 U161 ( .A1(\U6/DATA2_90 ), .A2(n626), .ZN(\U6/Z_90 ) );
  AND2_X1 U162 ( .A1(\U6/DATA2_9 ), .A2(n627), .ZN(\U6/Z_9 ) );
  AND2_X1 U163 ( .A1(\U6/DATA2_89 ), .A2(n627), .ZN(\U6/Z_89 ) );
  AND2_X1 U164 ( .A1(\U6/DATA2_88 ), .A2(n626), .ZN(\U6/Z_88 ) );
  AND2_X1 U165 ( .A1(\U6/DATA2_87 ), .A2(n627), .ZN(\U6/Z_87 ) );
  AND2_X1 U166 ( .A1(\U6/DATA2_86 ), .A2(n626), .ZN(\U6/Z_86 ) );
  AND2_X1 U167 ( .A1(\U6/DATA2_85 ), .A2(n627), .ZN(\U6/Z_85 ) );
  AND2_X1 U168 ( .A1(\U6/DATA2_84 ), .A2(n627), .ZN(\U6/Z_84 ) );
  AND2_X1 U169 ( .A1(\U6/DATA2_83 ), .A2(n626), .ZN(\U6/Z_83 ) );
  AND2_X1 U170 ( .A1(\U6/DATA2_82 ), .A2(n627), .ZN(\U6/Z_82 ) );
  AND2_X1 U171 ( .A1(\U6/DATA2_81 ), .A2(n627), .ZN(\U6/Z_81 ) );
  AND2_X1 U172 ( .A1(\U6/DATA2_80 ), .A2(n626), .ZN(\U6/Z_80 ) );
  AND2_X1 U173 ( .A1(\U6/DATA2_8 ), .A2(n626), .ZN(\U6/Z_8 ) );
  AND2_X1 U174 ( .A1(\U6/DATA2_79 ), .A2(n626), .ZN(\U6/Z_79 ) );
  AND2_X1 U175 ( .A1(\U6/DATA2_78 ), .A2(n627), .ZN(\U6/Z_78 ) );
  AND2_X1 U176 ( .A1(\U6/DATA2_77 ), .A2(n626), .ZN(\U6/Z_77 ) );
  AND2_X1 U177 ( .A1(\U6/DATA2_76 ), .A2(n627), .ZN(\U6/Z_76 ) );
  AND2_X1 U178 ( .A1(\U6/DATA2_75 ), .A2(n626), .ZN(\U6/Z_75 ) );
  AND2_X1 U179 ( .A1(\U6/DATA2_74 ), .A2(n627), .ZN(\U6/Z_74 ) );
  AND2_X1 U180 ( .A1(\U6/DATA2_73 ), .A2(n626), .ZN(\U6/Z_73 ) );
  AND2_X1 U181 ( .A1(\U6/DATA2_72 ), .A2(n626), .ZN(\U6/Z_72 ) );
  AND2_X1 U182 ( .A1(\U6/DATA2_71 ), .A2(n626), .ZN(\U6/Z_71 ) );
  AND2_X1 U183 ( .A1(\U6/DATA2_70 ), .A2(n627), .ZN(\U6/Z_70 ) );
  AND2_X1 U184 ( .A1(\U6/DATA2_7 ), .A2(n627), .ZN(\U6/Z_7 ) );
  AND2_X1 U185 ( .A1(\U6/DATA2_69 ), .A2(n626), .ZN(\U6/Z_69 ) );
  AND2_X1 U186 ( .A1(\U6/DATA2_68 ), .A2(n626), .ZN(\U6/Z_68 ) );
  AND2_X1 U187 ( .A1(\U6/DATA2_67 ), .A2(n627), .ZN(\U6/Z_67 ) );
  AND2_X1 U188 ( .A1(\U6/DATA2_66 ), .A2(n626), .ZN(\U6/Z_66 ) );
  AND2_X1 U189 ( .A1(\U6/DATA2_65 ), .A2(n627), .ZN(\U6/Z_65 ) );
  AND2_X1 U190 ( .A1(\U6/DATA2_64 ), .A2(n626), .ZN(\U6/Z_64 ) );
  AND2_X1 U191 ( .A1(\U6/DATA2_63 ), .A2(n627), .ZN(\U6/Z_63 ) );
  AND2_X1 U192 ( .A1(\U6/DATA2_62 ), .A2(n626), .ZN(\U6/Z_62 ) );
  AND2_X1 U193 ( .A1(\U6/DATA2_61 ), .A2(n627), .ZN(\U6/Z_61 ) );
  AND2_X1 U194 ( .A1(\U6/DATA2_60 ), .A2(n626), .ZN(\U6/Z_60 ) );
  AND2_X1 U195 ( .A1(\U6/DATA2_6 ), .A2(n627), .ZN(\U6/Z_6 ) );
  AND2_X1 U196 ( .A1(\U6/DATA2_59 ), .A2(n627), .ZN(\U6/Z_59 ) );
  AND2_X1 U197 ( .A1(\U6/DATA2_58 ), .A2(n626), .ZN(\U6/Z_58 ) );
  AND2_X1 U198 ( .A1(\U6/DATA2_57 ), .A2(n626), .ZN(\U6/Z_57 ) );
  AND2_X1 U199 ( .A1(\U6/DATA2_56 ), .A2(n626), .ZN(\U6/Z_56 ) );
  AND2_X1 U200 ( .A1(\U6/DATA2_55 ), .A2(n626), .ZN(\U6/Z_55 ) );
  AND2_X1 U201 ( .A1(\U6/DATA2_54 ), .A2(n626), .ZN(\U6/Z_54 ) );
  AND2_X1 U202 ( .A1(\U6/DATA2_53 ), .A2(n627), .ZN(\U6/Z_53 ) );
  AND2_X1 U203 ( .A1(\U6/DATA2_52 ), .A2(n627), .ZN(\U6/Z_52 ) );
  AND2_X1 U204 ( .A1(\U6/DATA2_51 ), .A2(n627), .ZN(\U6/Z_51 ) );
  AND2_X1 U205 ( .A1(\U6/DATA2_50 ), .A2(n627), .ZN(\U6/Z_50 ) );
  AND2_X1 U206 ( .A1(\U6/DATA2_5 ), .A2(n626), .ZN(\U6/Z_5 ) );
  AND2_X1 U207 ( .A1(\U6/DATA2_49 ), .A2(n626), .ZN(\U6/Z_49 ) );
  AND2_X1 U208 ( .A1(\U6/DATA2_48 ), .A2(n626), .ZN(\U6/Z_48 ) );
  AND2_X1 U209 ( .A1(\U6/DATA2_47 ), .A2(n627), .ZN(\U6/Z_47 ) );
  AND2_X1 U210 ( .A1(\U6/DATA2_46 ), .A2(n626), .ZN(\U6/Z_46 ) );
  AND2_X1 U211 ( .A1(\U6/DATA2_45 ), .A2(n627), .ZN(\U6/Z_45 ) );
  AND2_X1 U212 ( .A1(\U6/DATA2_44 ), .A2(n627), .ZN(\U6/Z_44 ) );
  AND2_X1 U213 ( .A1(\U6/DATA2_43 ), .A2(n627), .ZN(\U6/Z_43 ) );
  AND2_X1 U214 ( .A1(\U6/DATA2_42 ), .A2(n626), .ZN(\U6/Z_42 ) );
  AND2_X1 U215 ( .A1(\U6/DATA2_41 ), .A2(n627), .ZN(\U6/Z_41 ) );
  AND2_X1 U216 ( .A1(\U6/DATA2_40 ), .A2(n626), .ZN(\U6/Z_40 ) );
  AND2_X1 U217 ( .A1(\U6/DATA2_4 ), .A2(n627), .ZN(\U6/Z_4 ) );
  AND2_X1 U218 ( .A1(\U6/DATA2_39 ), .A2(n626), .ZN(\U6/Z_39 ) );
  AND2_X1 U219 ( .A1(\U6/DATA2_38 ), .A2(n627), .ZN(\U6/Z_38 ) );
  AND2_X1 U220 ( .A1(\U6/DATA2_37 ), .A2(n627), .ZN(\U6/Z_37 ) );
  AND2_X1 U221 ( .A1(\U6/DATA2_36 ), .A2(n626), .ZN(\U6/Z_36 ) );
  AND2_X1 U222 ( .A1(\U6/DATA2_35 ), .A2(n626), .ZN(\U6/Z_35 ) );
  AND2_X1 U223 ( .A1(\U6/DATA2_34 ), .A2(n627), .ZN(\U6/Z_34 ) );
  AND2_X1 U224 ( .A1(\U6/DATA2_33 ), .A2(n626), .ZN(\U6/Z_33 ) );
  AND2_X1 U225 ( .A1(\U6/DATA2_32 ), .A2(n627), .ZN(\U6/Z_32 ) );
  AND2_X1 U226 ( .A1(\U6/DATA2_31 ), .A2(n627), .ZN(\U6/Z_31 ) );
  AND2_X1 U227 ( .A1(\U6/DATA2_30 ), .A2(n626), .ZN(\U6/Z_30 ) );
  AND2_X1 U228 ( .A1(\U6/DATA2_3 ), .A2(n626), .ZN(\U6/Z_3 ) );
  AND2_X1 U229 ( .A1(\U6/DATA2_29 ), .A2(n627), .ZN(\U6/Z_29 ) );
  AND2_X1 U230 ( .A1(\U6/DATA2_28 ), .A2(n626), .ZN(\U6/Z_28 ) );
  AND2_X1 U231 ( .A1(\U6/DATA2_27 ), .A2(n626), .ZN(\U6/Z_27 ) );
  AND2_X1 U232 ( .A1(\U6/DATA2_26 ), .A2(n626), .ZN(\U6/Z_26 ) );
  AND2_X1 U233 ( .A1(\U6/DATA2_25 ), .A2(n626), .ZN(\U6/Z_25 ) );
  AND2_X1 U234 ( .A1(\U6/DATA2_24 ), .A2(n626), .ZN(\U6/Z_24 ) );
  AND2_X1 U235 ( .A1(\U6/DATA2_23 ), .A2(n626), .ZN(\U6/Z_23 ) );
  AND2_X1 U236 ( .A1(\U6/DATA2_22 ), .A2(n626), .ZN(\U6/Z_22 ) );
  AND2_X1 U237 ( .A1(\U6/DATA2_21 ), .A2(n626), .ZN(\U6/Z_21 ) );
  AND2_X1 U238 ( .A1(\U6/DATA2_20 ), .A2(n626), .ZN(\U6/Z_20 ) );
  AND2_X1 U239 ( .A1(\U6/DATA2_2 ), .A2(n626), .ZN(\U6/Z_2 ) );
  AND2_X1 U240 ( .A1(\U6/DATA2_19 ), .A2(n626), .ZN(\U6/Z_19 ) );
  AND2_X1 U241 ( .A1(\U6/DATA2_18 ), .A2(n626), .ZN(\U6/Z_18 ) );
  AND2_X1 U242 ( .A1(\U6/DATA2_17 ), .A2(n626), .ZN(\U6/Z_17 ) );
  AND2_X1 U243 ( .A1(\U6/DATA2_16 ), .A2(n627), .ZN(\U6/Z_16 ) );
  AND2_X1 U244 ( .A1(\U6/DATA2_15 ), .A2(n627), .ZN(\U6/Z_15 ) );
  AND2_X1 U245 ( .A1(\U6/DATA2_14 ), .A2(n627), .ZN(\U6/Z_14 ) );
  AND2_X1 U246 ( .A1(\U6/DATA2_13 ), .A2(n627), .ZN(\U6/Z_13 ) );
  AND2_X1 U247 ( .A1(\U6/DATA2_127 ), .A2(n627), .ZN(\U6/Z_127 ) );
  AND2_X1 U248 ( .A1(\U6/DATA2_126 ), .A2(n627), .ZN(\U6/Z_126 ) );
  AND2_X1 U249 ( .A1(\U6/DATA2_125 ), .A2(n627), .ZN(\U6/Z_125 ) );
  AND2_X1 U250 ( .A1(\U6/DATA2_124 ), .A2(n627), .ZN(\U6/Z_124 ) );
  AND2_X1 U251 ( .A1(\U6/DATA2_123 ), .A2(n627), .ZN(\U6/Z_123 ) );
  AND2_X1 U252 ( .A1(\U6/DATA2_122 ), .A2(n627), .ZN(\U6/Z_122 ) );
  AND2_X1 U253 ( .A1(\U6/DATA2_121 ), .A2(n627), .ZN(\U6/Z_121 ) );
  AND2_X1 U254 ( .A1(\U6/DATA2_120 ), .A2(n627), .ZN(\U6/Z_120 ) );
  AND2_X1 U255 ( .A1(\U6/DATA2_12 ), .A2(n627), .ZN(\U6/Z_12 ) );
  AND2_X1 U256 ( .A1(\U6/DATA2_119 ), .A2(n627), .ZN(\U6/Z_119 ) );
  AND2_X1 U257 ( .A1(\U6/DATA2_118 ), .A2(n626), .ZN(\U6/Z_118 ) );
  AND2_X1 U258 ( .A1(\U6/DATA2_117 ), .A2(n627), .ZN(\U6/Z_117 ) );
  AND2_X1 U259 ( .A1(\U6/DATA2_116 ), .A2(n626), .ZN(\U6/Z_116 ) );
  AND2_X1 U260 ( .A1(\U6/DATA2_115 ), .A2(n627), .ZN(\U6/Z_115 ) );
  AND2_X1 U261 ( .A1(\U6/DATA2_114 ), .A2(n626), .ZN(\U6/Z_114 ) );
  AND2_X1 U262 ( .A1(\U6/DATA2_113 ), .A2(n627), .ZN(\U6/Z_113 ) );
  AND2_X1 U263 ( .A1(\U6/DATA2_112 ), .A2(n626), .ZN(\U6/Z_112 ) );
  AND2_X1 U264 ( .A1(\U6/DATA2_111 ), .A2(n627), .ZN(\U6/Z_111 ) );
  AND2_X1 U265 ( .A1(\U6/DATA2_110 ), .A2(n626), .ZN(\U6/Z_110 ) );
  AND2_X1 U266 ( .A1(\U6/DATA2_11 ), .A2(n627), .ZN(\U6/Z_11 ) );
  AND2_X1 U267 ( .A1(\U6/DATA2_109 ), .A2(n626), .ZN(\U6/Z_109 ) );
  AND2_X1 U268 ( .A1(\U6/DATA2_108 ), .A2(n627), .ZN(\U6/Z_108 ) );
  AND2_X1 U269 ( .A1(\U6/DATA2_107 ), .A2(n627), .ZN(\U6/Z_107 ) );
  AND2_X1 U270 ( .A1(\U6/DATA2_106 ), .A2(n627), .ZN(\U6/Z_106 ) );
  AND2_X1 U271 ( .A1(\U6/DATA2_105 ), .A2(n626), .ZN(\U6/Z_105 ) );
  AND2_X1 U272 ( .A1(\U6/DATA2_104 ), .A2(n626), .ZN(\U6/Z_104 ) );
  AND2_X1 U273 ( .A1(\U6/DATA2_103 ), .A2(n626), .ZN(\U6/Z_103 ) );
  AND2_X1 U274 ( .A1(\U6/DATA2_102 ), .A2(n626), .ZN(\U6/Z_102 ) );
  AND2_X1 U275 ( .A1(\U6/DATA2_101 ), .A2(n626), .ZN(\U6/Z_101 ) );
  AND2_X1 U276 ( .A1(\U6/DATA2_100 ), .A2(n627), .ZN(\U6/Z_100 ) );
  AND2_X1 U277 ( .A1(\U6/DATA2_10 ), .A2(n627), .ZN(\U6/Z_10 ) );
  AND2_X1 U278 ( .A1(\U6/DATA2_1 ), .A2(n626), .ZN(\U6/Z_1 ) );
  AND2_X1 U279 ( .A1(\U6/DATA2_0 ), .A2(n626), .ZN(\U6/Z_0 ) );
  AND2_X1 U288 ( .A1(n142), .A2(n143), .ZN(n58) );
  AND2_X1 U289 ( .A1(n144), .A2(n142), .ZN(n57) );
  AND2_X1 U290 ( .A1(n720), .A2(n143), .ZN(n60) );
  AND2_X1 U291 ( .A1(n144), .A2(n720), .ZN(n59) );
  AND2_X1 U292 ( .A1(n624), .A2(n143), .ZN(n62) );
  AND2_X1 U293 ( .A1(n144), .A2(n624), .ZN(n61) );
  AND2_X1 U294 ( .A1(n144), .A2(n147), .ZN(n63) );
  AND2_X1 U295 ( .A1(n625), .A2(n142), .ZN(n70) );
  AND2_X1 U296 ( .A1(n142), .A2(n153), .ZN(n69) );
  AND2_X1 U297 ( .A1(n720), .A2(n625), .ZN(n72) );
  AND2_X1 U298 ( .A1(n720), .A2(n153), .ZN(n71) );
  AND2_X1 U299 ( .A1(n624), .A2(n625), .ZN(n74) );
  AND2_X1 U300 ( .A1(n624), .A2(n153), .ZN(n73) );
  AND2_X1 U301 ( .A1(n153), .A2(n147), .ZN(n75) );
  AND2_X1 U303 ( .A1(\U18/DATA1_0 ), .A2(start), .ZN(\U18/Z_0 ) );
  AND2_X1 U304 ( .A1(\U17/DATA1_0 ), .A2(start), .ZN(\U17/Z_0 ) );
  AND2_X1 U305 ( .A1(\U16/DATA1_0 ), .A2(start), .ZN(\U16/Z_0 ) );
  AND2_X1 U306 ( .A1(\U15/DATA1_0 ), .A2(start), .ZN(\U15/Z_0 ) );
  AND2_X1 U307 ( .A1(\U14/DATA1_0 ), .A2(start), .ZN(\U14/Z_0 ) );
  AND2_X1 U308 ( .A1(\U13/DATA1_0 ), .A2(start), .ZN(\U13/Z_0 ) );
  AND2_X1 U309 ( .A1(\U12/DATA1_0 ), .A2(start), .ZN(\U12/Z_0 ) );
  AND2_X1 U310 ( .A1(\U11/DATA1_0 ), .A2(start), .ZN(\U11/Z_0 ) );
  AND2_X1 U311 ( .A1(\U10/DATA1_0 ), .A2(start), .ZN(\U10/Z_0 ) );
  DFFR_X2 \ReadAddress_reg[0]  ( .D(n161), .CK(clock), .RN(n628), .Q(
        \add_101/A[0] ), .QN(n22) );
  DFF_X2 base_offset_reg ( .D(\U3/U1/DATA2_15 ), .CK(clock), .Q(DataOut[15])
         );
  DFFR_X2 \ReadAddress_reg[2]  ( .D(n723), .CK(clock), .RN(n628), .Q(
        \add_101/A[2] ), .QN(n650) );
  DFFR_X2 \ReadAddress_reg[12]  ( .D(n733), .CK(clock), .RN(n629), .Q(
        \add_101/A[12] ), .QN(n694) );
  DFFR_X2 \ReadAddress_reg[10]  ( .D(n731), .CK(clock), .RN(n629), .Q(
        \add_101/A[10] ), .QN(n685) );
  DFFR_X2 \ReadAddress_reg[8]  ( .D(n729), .CK(clock), .RN(n628), .Q(
        \add_101/A[8] ), .QN(n676) );
  DFFR_X2 \ReadAddress_reg[6]  ( .D(n727), .CK(clock), .RN(n628), .Q(
        \add_101/A[6] ), .QN(n667) );
  DFFR_X2 \ReadAddress_reg[4]  ( .D(n725), .CK(clock), .RN(n628), .Q(
        \add_101/A[4] ), .QN(n658) );
  DFFR_X2 \ReadAddress_reg[13]  ( .D(n734), .CK(clock), .RN(n629), .Q(
        \add_101/A[13] ), .QN(n698) );
  DFFR_X2 \ReadAddress_reg[1]  ( .D(n722), .CK(clock), .RN(n628), .Q(
        \add_101/A[1] ) );
  DFFR_X2 \ReadAddress_reg[11]  ( .D(n732), .CK(clock), .RN(n629), .Q(
        \add_101/A[11] ), .QN(n642) );
  DFFR_X2 \ReadAddress_reg[9]  ( .D(n730), .CK(clock), .RN(n629), .Q(
        \add_101/A[9] ), .QN(n641) );
  DFFR_X2 \ReadAddress_reg[7]  ( .D(n728), .CK(clock), .RN(n628), .Q(
        \add_101/A[7] ) );
  DFFR_X2 \ReadAddress_reg[5]  ( .D(n726), .CK(clock), .RN(n628), .Q(
        \add_101/A[5] ) );
  DFFR_X2 \ReadAddress_reg[3]  ( .D(n724), .CK(clock), .RN(n628), .Q(
        \add_101/A[3] ) );
  DFFR_X2 \ReadAddress_reg[14]  ( .D(n735), .CK(clock), .RN(n629), .Q(
        \add_101/A[14] ), .QN(n708) );
  DFFR_X2 \ReadAddress_reg[15]  ( .D(n736), .CK(clock), .RN(n629), .Q(
        \add_101/A[15] ) );
  INV_X4 U4 ( .A(1'b1), .ZN(DataOut[8]) );
  INV_X4 U6 ( .A(1'b1), .ZN(DataOut[9]) );
  INV_X4 U8 ( .A(1'b1), .ZN(DataOut[10]) );
  INV_X4 U10 ( .A(1'b1), .ZN(DataOut[11]) );
  INV_X4 U12 ( .A(1'b1), .ZN(DataOut[12]) );
  INV_X4 U14 ( .A(1'b1), .ZN(DataOut[13]) );
  INV_X4 U16 ( .A(1'b1), .ZN(DataOut[14]) );
  AND2_X4 U18 ( .A1(n48), .A2(n737), .ZN(n623) );
  AND2_X4 U19 ( .A1(n26), .A2(\add_95/A[2] ), .ZN(n624) );
  AND2_X4 U20 ( .A1(n24), .A2(\add_95/A[0] ), .ZN(n625) );
  NAND2_X1 U21 ( .A1(\U3/U1/DATA2_15 ), .A2(n709), .ZN(n716) );
  OR2_X4 U22 ( .A1(n51), .A2(n52), .ZN(\U5/Z_7 ) );
  OR2_X4 U23 ( .A1(n76), .A2(n77), .ZN(\U5/Z_6 ) );
  OR2_X4 U24 ( .A1(n86), .A2(n87), .ZN(\U5/Z_5 ) );
  OR2_X4 U26 ( .A1(n96), .A2(n97), .ZN(\U5/Z_4 ) );
  OR2_X4 U27 ( .A1(n106), .A2(n107), .ZN(\U5/Z_3 ) );
  OR2_X4 U28 ( .A1(n116), .A2(n117), .ZN(\U5/Z_2 ) );
  OR2_X4 U29 ( .A1(n126), .A2(n127), .ZN(\U5/Z_1 ) );
  OR2_X4 U31 ( .A1(n136), .A2(n137), .ZN(\U5/Z_0 ) );
  NAND2_X1 U32 ( .A1(\add_101/A[13] ), .A2(n701), .ZN(n707) );
  NOR4_X1 U33 ( .A1(\add_101/A[12] ), .A2(\add_101/A[10] ), .A3(
        \add_101/A[13] ), .A4(n709), .ZN(n645) );
  XOR2_X1 U34 ( .A(n700), .B(\add_101/A[13] ), .Z(n699) );
  INV_X4 U36 ( .A(n639), .ZN(n631) );
  INV_X4 U37 ( .A(n639), .ZN(n630) );
  INV_X4 U38 ( .A(n639), .ZN(n632) );
  INV_X4 U39 ( .A(n639), .ZN(n636) );
  INV_X4 U41 ( .A(n639), .ZN(n635) );
  INV_X4 U42 ( .A(n639), .ZN(n634) );
  INV_X4 U43 ( .A(n639), .ZN(n633) );
  INV_X4 U44 ( .A(n639), .ZN(n629) );
  INV_X4 U46 ( .A(n639), .ZN(n628) );
  INV_X4 U47 ( .A(n639), .ZN(n637) );
  INV_X4 U48 ( .A(n623), .ZN(n626) );
  INV_X4 U49 ( .A(n623), .ZN(n627) );
  INV_X4 U51 ( .A(n639), .ZN(n638) );
  INV_X4 U52 ( .A(reset_n), .ZN(n639) );
  AOI22_X2 U53 ( .A1(\U5/DATA10_0 ), .A2(n75), .B1(\U5/DATA9_0 ), .B2(n738), 
        .ZN(n148) );
  AOI22_X2 U54 ( .A1(\U5/DATA10_1 ), .A2(n75), .B1(\U5/DATA9_1 ), .B2(n738), 
        .ZN(n132) );
  AOI22_X2 U56 ( .A1(\U5/DATA10_2 ), .A2(n75), .B1(\U5/DATA9_2 ), .B2(n738), 
        .ZN(n122) );
  AOI22_X2 U57 ( .A1(\U5/DATA10_3 ), .A2(n75), .B1(\U5/DATA9_3 ), .B2(n738), 
        .ZN(n112) );
  AOI22_X2 U58 ( .A1(\U5/DATA10_4 ), .A2(n75), .B1(\U5/DATA9_4 ), .B2(n738), 
        .ZN(n102) );
  AOI22_X2 U59 ( .A1(\U5/DATA10_5 ), .A2(n75), .B1(\U5/DATA9_5 ), .B2(n738), 
        .ZN(n92) );
  AOI22_X1 U61 ( .A1(\U5/DATA10_6 ), .A2(n75), .B1(\U5/DATA9_6 ), .B2(n738), 
        .ZN(n82) );
  AOI22_X1 U62 ( .A1(\U5/DATA10_7 ), .A2(n75), .B1(\U5/DATA9_7 ), .B2(n738), 
        .ZN(n65) );
  NAND2_X2 U63 ( .A1(n704), .A2(start), .ZN(n737) );
  AOI22_X2 U64 ( .A1(\U5/DATA2_0 ), .A2(n63), .B1(\U5/DATA1_0 ), .B2(n64), 
        .ZN(n138) );
  AOI22_X2 U66 ( .A1(\U5/DATA2_1 ), .A2(n63), .B1(\U5/DATA1_1 ), .B2(n64), 
        .ZN(n128) );
  AOI22_X2 U67 ( .A1(\U5/DATA2_2 ), .A2(n63), .B1(\U5/DATA1_2 ), .B2(n64), 
        .ZN(n118) );
  AOI22_X2 U68 ( .A1(\U5/DATA2_3 ), .A2(n63), .B1(\U5/DATA1_3 ), .B2(n64), 
        .ZN(n108) );
  AOI22_X2 U69 ( .A1(\U5/DATA2_4 ), .A2(n63), .B1(\U5/DATA1_4 ), .B2(n64), 
        .ZN(n98) );
  AOI22_X2 U71 ( .A1(\U5/DATA2_5 ), .A2(n63), .B1(\U5/DATA1_5 ), .B2(n64), 
        .ZN(n88) );
  AOI22_X1 U72 ( .A1(\U5/DATA2_6 ), .A2(n63), .B1(\U5/DATA1_6 ), .B2(n64), 
        .ZN(n78) );
  AOI22_X1 U73 ( .A1(\U5/DATA2_7 ), .A2(n63), .B1(\U5/DATA1_7 ), .B2(n64), 
        .ZN(n53) );
  AOI22_X2 U74 ( .A1(\U5/DATA4_0 ), .A2(n61), .B1(\U5/DATA3_0 ), .B2(n62), 
        .ZN(n139) );
  AOI22_X2 U76 ( .A1(\U5/DATA12_0 ), .A2(n73), .B1(\U5/DATA11_0 ), .B2(n74), 
        .ZN(n149) );
  AOI22_X2 U77 ( .A1(\U5/DATA4_1 ), .A2(n61), .B1(\U5/DATA3_1 ), .B2(n62), 
        .ZN(n129) );
  AOI22_X2 U78 ( .A1(\U5/DATA12_1 ), .A2(n73), .B1(\U5/DATA11_1 ), .B2(n74), 
        .ZN(n133) );
  AOI22_X2 U79 ( .A1(\U5/DATA4_2 ), .A2(n61), .B1(\U5/DATA3_2 ), .B2(n62), 
        .ZN(n119) );
  AOI22_X2 U81 ( .A1(\U5/DATA12_2 ), .A2(n73), .B1(\U5/DATA11_2 ), .B2(n74), 
        .ZN(n123) );
  AOI22_X2 U82 ( .A1(\U5/DATA4_3 ), .A2(n61), .B1(\U5/DATA3_3 ), .B2(n62), 
        .ZN(n109) );
  AOI22_X2 U83 ( .A1(\U5/DATA12_3 ), .A2(n73), .B1(\U5/DATA11_3 ), .B2(n74), 
        .ZN(n113) );
  AOI22_X2 U84 ( .A1(\U5/DATA4_4 ), .A2(n61), .B1(\U5/DATA3_4 ), .B2(n62), 
        .ZN(n99) );
  AOI22_X2 U86 ( .A1(\U5/DATA12_4 ), .A2(n73), .B1(\U5/DATA11_4 ), .B2(n74), 
        .ZN(n103) );
  AOI22_X2 U87 ( .A1(\U5/DATA4_5 ), .A2(n61), .B1(\U5/DATA3_5 ), .B2(n62), 
        .ZN(n89) );
  AOI22_X2 U88 ( .A1(\U5/DATA12_5 ), .A2(n73), .B1(\U5/DATA11_5 ), .B2(n74), 
        .ZN(n93) );
  AOI22_X1 U89 ( .A1(\U5/DATA4_6 ), .A2(n61), .B1(\U5/DATA3_6 ), .B2(n62), 
        .ZN(n79) );
  AOI22_X1 U91 ( .A1(\U5/DATA12_6 ), .A2(n73), .B1(\U5/DATA11_6 ), .B2(n74), 
        .ZN(n83) );
  AOI22_X1 U92 ( .A1(\U5/DATA4_7 ), .A2(n61), .B1(\U5/DATA3_7 ), .B2(n62), 
        .ZN(n54) );
  AOI22_X1 U93 ( .A1(\U5/DATA12_7 ), .A2(n73), .B1(\U5/DATA11_7 ), .B2(n74), 
        .ZN(n66) );
  AOI22_X2 U94 ( .A1(\U5/DATA8_0 ), .A2(n57), .B1(\U5/DATA7_0 ), .B2(n58), 
        .ZN(n141) );
  AOI22_X2 U96 ( .A1(\U5/DATA6_0 ), .A2(n59), .B1(\U5/DATA5_0 ), .B2(n60), 
        .ZN(n140) );
  AOI22_X2 U97 ( .A1(\U5/DATA16_0 ), .A2(n69), .B1(\U5/DATA15_0 ), .B2(n70), 
        .ZN(n151) );
  AOI22_X2 U98 ( .A1(\U5/DATA14_0 ), .A2(n71), .B1(\U5/DATA13_0 ), .B2(n72), 
        .ZN(n150) );
  AOI22_X2 U99 ( .A1(\U5/DATA8_1 ), .A2(n57), .B1(\U5/DATA7_1 ), .B2(n58), 
        .ZN(n131) );
  AOI22_X2 U102 ( .A1(\U5/DATA6_1 ), .A2(n59), .B1(\U5/DATA5_1 ), .B2(n60), 
        .ZN(n130) );
  AOI22_X2 U104 ( .A1(\U5/DATA16_1 ), .A2(n69), .B1(\U5/DATA15_1 ), .B2(n70), 
        .ZN(n135) );
  AOI22_X2 U105 ( .A1(\U5/DATA14_1 ), .A2(n71), .B1(\U5/DATA13_1 ), .B2(n72), 
        .ZN(n134) );
  AOI22_X2 U106 ( .A1(\U5/DATA8_2 ), .A2(n57), .B1(\U5/DATA7_2 ), .B2(n58), 
        .ZN(n121) );
  AOI22_X2 U110 ( .A1(\U5/DATA6_2 ), .A2(n59), .B1(\U5/DATA5_2 ), .B2(n60), 
        .ZN(n120) );
  AOI22_X2 U112 ( .A1(\U5/DATA16_2 ), .A2(n69), .B1(\U5/DATA15_2 ), .B2(n70), 
        .ZN(n125) );
  AOI22_X2 U113 ( .A1(\U5/DATA14_2 ), .A2(n71), .B1(\U5/DATA13_2 ), .B2(n72), 
        .ZN(n124) );
  AOI22_X2 U114 ( .A1(\U5/DATA8_3 ), .A2(n57), .B1(\U5/DATA7_3 ), .B2(n58), 
        .ZN(n111) );
  AOI22_X2 U119 ( .A1(\U5/DATA6_3 ), .A2(n59), .B1(\U5/DATA5_3 ), .B2(n60), 
        .ZN(n110) );
  AOI22_X2 U120 ( .A1(\U5/DATA16_3 ), .A2(n69), .B1(\U5/DATA15_3 ), .B2(n70), 
        .ZN(n115) );
  AOI22_X2 U121 ( .A1(\U5/DATA14_3 ), .A2(n71), .B1(\U5/DATA13_3 ), .B2(n72), 
        .ZN(n114) );
  AOI22_X2 U122 ( .A1(\U5/DATA8_4 ), .A2(n57), .B1(\U5/DATA7_4 ), .B2(n58), 
        .ZN(n101) );
  AOI22_X2 U123 ( .A1(\U5/DATA6_4 ), .A2(n59), .B1(\U5/DATA5_4 ), .B2(n60), 
        .ZN(n100) );
  AOI22_X2 U124 ( .A1(\U5/DATA16_4 ), .A2(n69), .B1(\U5/DATA15_4 ), .B2(n70), 
        .ZN(n105) );
  AOI22_X2 U127 ( .A1(\U5/DATA14_4 ), .A2(n71), .B1(\U5/DATA13_4 ), .B2(n72), 
        .ZN(n104) );
  AOI22_X2 U128 ( .A1(\U5/DATA8_5 ), .A2(n57), .B1(\U5/DATA7_5 ), .B2(n58), 
        .ZN(n91) );
  AOI22_X2 U129 ( .A1(\U5/DATA6_5 ), .A2(n59), .B1(\U5/DATA5_5 ), .B2(n60), 
        .ZN(n90) );
  AOI22_X2 U130 ( .A1(\U5/DATA16_5 ), .A2(n69), .B1(\U5/DATA15_5 ), .B2(n70), 
        .ZN(n95) );
  AOI22_X2 U131 ( .A1(\U5/DATA14_5 ), .A2(n71), .B1(\U5/DATA13_5 ), .B2(n72), 
        .ZN(n94) );
  AOI22_X1 U132 ( .A1(\U5/DATA8_6 ), .A2(n57), .B1(\U5/DATA7_6 ), .B2(n58), 
        .ZN(n81) );
  AOI22_X1 U133 ( .A1(\U5/DATA6_6 ), .A2(n59), .B1(\U5/DATA5_6 ), .B2(n60), 
        .ZN(n80) );
  AOI22_X1 U134 ( .A1(\U5/DATA16_6 ), .A2(n69), .B1(\U5/DATA15_6 ), .B2(n70), 
        .ZN(n85) );
  AOI22_X1 U135 ( .A1(\U5/DATA14_6 ), .A2(n71), .B1(\U5/DATA13_6 ), .B2(n72), 
        .ZN(n84) );
  AOI22_X1 U136 ( .A1(\U5/DATA8_7 ), .A2(n57), .B1(\U5/DATA7_7 ), .B2(n58), 
        .ZN(n56) );
  AOI22_X1 U137 ( .A1(\U5/DATA6_7 ), .A2(n59), .B1(\U5/DATA5_7 ), .B2(n60), 
        .ZN(n55) );
  AOI22_X1 U138 ( .A1(\U5/DATA16_7 ), .A2(n69), .B1(\U5/DATA15_7 ), .B2(n70), 
        .ZN(n68) );
  AOI22_X1 U139 ( .A1(\U5/DATA14_7 ), .A2(n71), .B1(\U5/DATA13_7 ), .B2(n72), 
        .ZN(n67) );
  OAI21_X2 U140 ( .B1(n22), .B2(n704), .A(n703), .ZN(n161) );
  AND2_X4 U141 ( .A1(n147), .A2(n143), .ZN(n64) );
  INV_X4 U142 ( .A(n64), .ZN(n640) );
  NAND2_X2 U143 ( .A1(start), .A2(n640), .ZN(n717) );
  NOR4_X2 U144 ( .A1(n642), .A2(n708), .A3(n676), .A4(n641), .ZN(n646) );
  INV_X4 U145 ( .A(start), .ZN(n709) );
  NOR4_X2 U146 ( .A1(\add_101/A[5] ), .A2(\add_101/A[4] ), .A3(\add_101/A[7] ), 
        .A4(\add_101/A[6] ), .ZN(n644) );
  NOR4_X2 U147 ( .A1(\add_101/A[1] ), .A2(\add_101/A[0] ), .A3(\add_101/A[3] ), 
        .A4(\add_101/A[2] ), .ZN(n643) );
  NAND4_X2 U148 ( .A1(n646), .A2(n645), .A3(n644), .A4(n643), .ZN(n50) );
  NAND2_X2 U280 ( .A1(n717), .A2(n50), .ZN(n711) );
  INV_X4 U281 ( .A(n711), .ZN(n704) );
  NOR2_X2 U282 ( .A1(n737), .A2(n22), .ZN(n647) );
  INV_X4 U283 ( .A(n737), .ZN(n706) );
  NAND2_X2 U284 ( .A1(n706), .A2(n22), .ZN(n703) );
  NAND2_X2 U285 ( .A1(n704), .A2(n703), .ZN(n649) );
  MUX2_X2 U286 ( .A(n647), .B(n649), .S(\add_101/A[1] ), .Z(n722) );
  NAND2_X2 U287 ( .A1(\add_101/A[0] ), .A2(n650), .ZN(n648) );
  MUX2_X2 U302 ( .A(n650), .B(n648), .S(\add_101/A[1] ), .Z(n652) );
  INV_X4 U312 ( .A(n649), .ZN(n651) );
  OAI22_X2 U313 ( .A1(n737), .A2(n652), .B1(n651), .B2(n650), .ZN(n723) );
  NAND3_X2 U314 ( .A1(\add_101/A[1] ), .A2(\add_101/A[0] ), .A3(\add_101/A[2] ), .ZN(n655) );
  NOR2_X2 U315 ( .A1(n737), .A2(n655), .ZN(n654) );
  NAND2_X2 U316 ( .A1(n655), .A2(n706), .ZN(n653) );
  NAND2_X2 U317 ( .A1(n704), .A2(n653), .ZN(n657) );
  MUX2_X2 U318 ( .A(n654), .B(n657), .S(\add_101/A[3] ), .Z(n724) );
  INV_X4 U319 ( .A(n655), .ZN(n661) );
  NAND2_X2 U320 ( .A1(n661), .A2(n658), .ZN(n656) );
  MUX2_X2 U321 ( .A(n658), .B(n656), .S(\add_101/A[3] ), .Z(n660) );
  INV_X4 U322 ( .A(n657), .ZN(n659) );
  OAI22_X2 U323 ( .A1(n737), .A2(n660), .B1(n659), .B2(n658), .ZN(n725) );
  NAND3_X2 U324 ( .A1(\add_101/A[4] ), .A2(\add_101/A[3] ), .A3(n661), .ZN(
        n664) );
  NOR2_X2 U325 ( .A1(n737), .A2(n664), .ZN(n663) );
  NAND2_X2 U326 ( .A1(n664), .A2(n706), .ZN(n662) );
  NAND2_X2 U327 ( .A1(n704), .A2(n662), .ZN(n666) );
  MUX2_X2 U328 ( .A(n663), .B(n666), .S(\add_101/A[5] ), .Z(n726) );
  INV_X4 U329 ( .A(n664), .ZN(n670) );
  NAND2_X2 U330 ( .A1(n670), .A2(n667), .ZN(n665) );
  MUX2_X2 U331 ( .A(n667), .B(n665), .S(\add_101/A[5] ), .Z(n669) );
  INV_X4 U332 ( .A(n666), .ZN(n668) );
  OAI22_X2 U333 ( .A1(n737), .A2(n669), .B1(n668), .B2(n667), .ZN(n727) );
  NAND3_X2 U334 ( .A1(\add_101/A[6] ), .A2(\add_101/A[5] ), .A3(n670), .ZN(
        n673) );
  NOR2_X2 U335 ( .A1(n737), .A2(n673), .ZN(n672) );
  NAND2_X2 U336 ( .A1(n673), .A2(n706), .ZN(n671) );
  NAND2_X2 U337 ( .A1(n704), .A2(n671), .ZN(n675) );
  MUX2_X2 U338 ( .A(n672), .B(n675), .S(\add_101/A[7] ), .Z(n728) );
  INV_X4 U339 ( .A(n673), .ZN(n679) );
  NAND2_X2 U340 ( .A1(n679), .A2(n676), .ZN(n674) );
  MUX2_X2 U341 ( .A(n676), .B(n674), .S(\add_101/A[7] ), .Z(n678) );
  INV_X4 U342 ( .A(n675), .ZN(n677) );
  OAI22_X2 U343 ( .A1(n737), .A2(n678), .B1(n677), .B2(n676), .ZN(n729) );
  NAND3_X2 U344 ( .A1(\add_101/A[7] ), .A2(\add_101/A[8] ), .A3(n679), .ZN(
        n682) );
  NOR2_X2 U345 ( .A1(n737), .A2(n682), .ZN(n681) );
  NAND2_X2 U346 ( .A1(n682), .A2(n706), .ZN(n680) );
  NAND2_X2 U347 ( .A1(n704), .A2(n680), .ZN(n684) );
  MUX2_X2 U348 ( .A(n681), .B(n684), .S(\add_101/A[9] ), .Z(n730) );
  INV_X4 U349 ( .A(n682), .ZN(n688) );
  NAND2_X2 U350 ( .A1(n688), .A2(n685), .ZN(n683) );
  MUX2_X2 U351 ( .A(n685), .B(n683), .S(\add_101/A[9] ), .Z(n687) );
  INV_X4 U352 ( .A(n684), .ZN(n686) );
  OAI22_X2 U353 ( .A1(n737), .A2(n687), .B1(n686), .B2(n685), .ZN(n731) );
  NAND3_X2 U354 ( .A1(\add_101/A[10] ), .A2(\add_101/A[9] ), .A3(n688), .ZN(
        n691) );
  NOR2_X2 U355 ( .A1(n737), .A2(n691), .ZN(n690) );
  NAND2_X2 U356 ( .A1(n691), .A2(n706), .ZN(n689) );
  NAND2_X2 U357 ( .A1(n704), .A2(n689), .ZN(n693) );
  MUX2_X2 U358 ( .A(n690), .B(n693), .S(\add_101/A[11] ), .Z(n732) );
  INV_X4 U359 ( .A(n691), .ZN(n697) );
  NAND2_X2 U360 ( .A1(n697), .A2(n694), .ZN(n692) );
  MUX2_X2 U361 ( .A(n694), .B(n692), .S(\add_101/A[11] ), .Z(n696) );
  INV_X4 U362 ( .A(n693), .ZN(n695) );
  OAI22_X2 U363 ( .A1(n737), .A2(n696), .B1(n695), .B2(n694), .ZN(n733) );
  NAND3_X2 U364 ( .A1(\add_101/A[12] ), .A2(\add_101/A[11] ), .A3(n697), .ZN(
        n700) );
  OAI22_X2 U365 ( .A1(n737), .A2(n699), .B1(n704), .B2(n698), .ZN(n734) );
  INV_X4 U366 ( .A(n700), .ZN(n701) );
  XOR2_X2 U367 ( .A(n707), .B(\add_101/A[14] ), .Z(n702) );
  OAI22_X2 U368 ( .A1(n737), .A2(n702), .B1(n704), .B2(n708), .ZN(n735) );
  INV_X4 U369 ( .A(n707), .ZN(n705) );
  NAND3_X2 U370 ( .A1(\add_101/A[14] ), .A2(n706), .A3(n705), .ZN(n714) );
  NOR2_X2 U371 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X2 U372 ( .A1(n710), .A2(n709), .ZN(n712) );
  NOR2_X2 U373 ( .A1(n712), .A2(n711), .ZN(n713) );
  MUX2_X2 U374 ( .A(n714), .B(n713), .S(\add_101/A[15] ), .Z(n715) );
  NAND2_X2 U375 ( .A1(n716), .A2(n715), .ZN(n736) );
  NAND2_X2 U376 ( .A1(\add_95/A[1] ), .A2(n25), .ZN(n718) );
  INV_X4 U377 ( .A(n718), .ZN(n720) );
  INV_X4 U378 ( .A(n717), .ZN(n49) );
  NOR2_X2 U379 ( .A1(n718), .A2(n27), .ZN(n719) );
  NOR2_X2 U380 ( .A1(n624), .A2(n719), .ZN(n155) );
  INV_X4 U381 ( .A(n50), .ZN(n739) );
  INV_X4 U382 ( .A(\U4/Z_0 ), .ZN(n721) );
  INV_X4 U383 ( .A(n154), .ZN(n738) );
endmodule


module Output_Fetch_Cdf ( clock, reset_n, ReadBus, DataOut, StartIn, StartOut
 );
  input [19:0] ReadBus;
  output [19:0] DataOut;
  input clock, reset_n, StartIn;
  output StartOut;
  wire   \U3/U1/Z_0 ;
  assign \U3/U1/Z_0  = StartIn;

  DFF_X1 \DataOut_reg[19]  ( .D(ReadBus[19]), .CK(clock), .Q(DataOut[19]) );
  DFF_X1 \DataOut_reg[18]  ( .D(ReadBus[18]), .CK(clock), .Q(DataOut[18]) );
  DFF_X1 \DataOut_reg[17]  ( .D(ReadBus[17]), .CK(clock), .Q(DataOut[17]) );
  DFF_X1 \DataOut_reg[16]  ( .D(ReadBus[16]), .CK(clock), .Q(DataOut[16]) );
  DFF_X1 \DataOut_reg[15]  ( .D(ReadBus[15]), .CK(clock), .Q(DataOut[15]) );
  DFF_X1 \DataOut_reg[14]  ( .D(ReadBus[14]), .CK(clock), .Q(DataOut[14]) );
  DFF_X1 \DataOut_reg[13]  ( .D(ReadBus[13]), .CK(clock), .Q(DataOut[13]) );
  DFF_X1 \DataOut_reg[12]  ( .D(ReadBus[12]), .CK(clock), .Q(DataOut[12]) );
  DFF_X1 \DataOut_reg[11]  ( .D(ReadBus[11]), .CK(clock), .Q(DataOut[11]) );
  DFF_X1 \DataOut_reg[10]  ( .D(ReadBus[10]), .CK(clock), .Q(DataOut[10]) );
  DFF_X1 \DataOut_reg[9]  ( .D(ReadBus[9]), .CK(clock), .Q(DataOut[9]) );
  DFF_X1 \DataOut_reg[8]  ( .D(ReadBus[8]), .CK(clock), .Q(DataOut[8]) );
  DFF_X1 \DataOut_reg[7]  ( .D(ReadBus[7]), .CK(clock), .Q(DataOut[7]) );
  DFF_X1 \DataOut_reg[6]  ( .D(ReadBus[6]), .CK(clock), .Q(DataOut[6]) );
  DFF_X1 \DataOut_reg[5]  ( .D(ReadBus[5]), .CK(clock), .Q(DataOut[5]) );
  DFF_X1 \DataOut_reg[4]  ( .D(ReadBus[4]), .CK(clock), .Q(DataOut[4]) );
  DFF_X1 \DataOut_reg[3]  ( .D(ReadBus[3]), .CK(clock), .Q(DataOut[3]) );
  DFF_X1 \DataOut_reg[2]  ( .D(ReadBus[2]), .CK(clock), .Q(DataOut[2]) );
  DFF_X1 \DataOut_reg[1]  ( .D(ReadBus[1]), .CK(clock), .Q(DataOut[1]) );
  DFF_X1 \DataOut_reg[0]  ( .D(ReadBus[0]), .CK(clock), .Q(DataOut[0]) );
  DFFR_X2 StartOut_reg ( .D(\U3/U1/Z_0 ), .CK(clock), .RN(reset_n), .Q(
        StartOut) );
endmodule


module Output_TopExpression ( clock, reset_n, DataIn, CdfMin, StartIn, 
        StartOut, DataOut );
  input [19:0] DataIn;
  input [19:0] CdfMin;
  output [27:0] DataOut;
  input clock, reset_n, StartIn;
  output StartOut;
  wire   n81, n162, \U8/Z_0 , \U8/Z_1 , \U8/Z_2 , \U8/Z_3 , \U8/Z_4 , \U8/Z_5 ,
         \U8/Z_6 , \U8/Z_7 , \U8/Z_8 , \U8/Z_9 , \U8/Z_10 , \U8/Z_11 ,
         \U8/Z_12 , \U8/Z_13 , \U8/DATA1_8 , \U8/DATA1_9 , \U8/DATA1_10 ,
         \U8/DATA1_11 , \U8/DATA1_12 , \U8/DATA1_13 , \U7/Z_1 , \U7/Z_2 ,
         \U7/Z_3 , \U7/Z_4 , \U7/Z_5 , \U7/Z_6 , \U7/Z_7 , \U7/Z_8 , \U7/Z_9 ,
         \U7/Z_10 , \U7/Z_11 , \U7/Z_12 , \U7/Z_13 , \U7/Z_14 , \U7/Z_15 ,
         \U7/Z_16 , \U7/Z_17 , \U7/Z_18 , \U7/Z_19 , \U7/DATA1_0 , \U6/Z_1 ,
         \U6/Z_2 , \U6/Z_3 , \U6/Z_4 , \U6/Z_5 , \U6/Z_6 , \U6/Z_7 , \U6/Z_8 ,
         \U6/Z_9 , \U6/Z_10 , \U6/Z_11 , \U6/Z_12 , \U6/Z_13 , \U5/Z_0 ,
         \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 ,
         \U4/Z_7 , \U4/Z_8 , \U4/Z_9 , \U4/Z_10 , \U4/Z_11 , \U4/Z_12 ,
         \U4/Z_13 , \U4/Z_14 , \U4/Z_15 , \U4/Z_16 , \U4/Z_17 , \U4/Z_18 ,
         \U4/Z_19 , \U4/Z_20 , \U4/Z_21 , \U4/Z_22 , \U4/Z_23 , \U4/Z_24 ,
         \U4/Z_25 , \U4/Z_26 , \U4/Z_27 , \U4/DATA1_0 , \U4/DATA1_1 ,
         \U4/DATA1_2 , \U4/DATA1_3 , \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 ,
         \U4/DATA1_7 , \U4/DATA1_8 , \U4/DATA1_9 , \U4/DATA1_10 ,
         \U4/DATA1_11 , \U4/DATA1_12 , \U4/DATA1_13 , \top_add/CI ,
         \top_add/A[0] , \top_add/A[1] , \top_add/A[2] , \top_add/A[3] ,
         \top_add/A[4] , \top_add/A[5] , \top_add/A[11] , \top_add/A[12] ,
         \top_add/A[13] , \bottom_add/A[8] , \bottom_add/A[9] ,
         \bottom_add/A[10] , \bottom_add/A[11] , \bottom_add/A[12] ,
         \bottom_add/A[13] , \first_add/A[0] , \first_add/A[1] ,
         \first_add/A[2] , \first_add/A[3] , \first_add/A[4] ,
         \first_add/A[5] , \first_add/A[6] , \first_add/A[7] ,
         \first_add/A[8] , \first_add/A[9] , \first_add/A[10] ,
         \first_add/A[11] , \first_add/A[12] , \first_add/A[13] ,
         \first_add/A[14] , \first_add/A[15] , \first_add/A[16] ,
         \first_add/A[17] , \first_add/A[18] , \first_add/A[19] , n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n20, n21, n22, n23,
         n24, n25, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603;
  assign \first_add/A[0]  = DataIn[0];
  assign \first_add/A[1]  = DataIn[1];
  assign \first_add/A[2]  = DataIn[2];
  assign \first_add/A[3]  = DataIn[3];
  assign \first_add/A[4]  = DataIn[4];
  assign \first_add/A[5]  = DataIn[5];
  assign \first_add/A[6]  = DataIn[6];
  assign \first_add/A[7]  = DataIn[7];
  assign \first_add/A[8]  = DataIn[8];
  assign \first_add/A[9]  = DataIn[9];
  assign \first_add/A[10]  = DataIn[10];
  assign \first_add/A[11]  = DataIn[11];
  assign \first_add/A[12]  = DataIn[12];
  assign \first_add/A[13]  = DataIn[13];
  assign \first_add/A[14]  = DataIn[14];
  assign \first_add/A[15]  = DataIn[15];
  assign \first_add/A[16]  = DataIn[16];
  assign \first_add/A[17]  = DataIn[17];
  assign \first_add/A[18]  = DataIn[18];
  assign \first_add/A[19]  = DataIn[19];

  DFFR_X1 \Data_reg[5]  ( .D(\U7/Z_5 ), .CK(clock), .RN(n339), .Q(
        \bottom_add/A[13] ), .QN(n14) );
  DFFR_X1 \Data_reg[4]  ( .D(\U7/Z_4 ), .CK(clock), .RN(n339), .Q(
        \bottom_add/A[12] ), .QN(n15) );
  DFFR_X1 \Data_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .RN(n339), .Q(
        \bottom_add/A[11] ), .QN(n16) );
  DFFR_X1 \Data_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .RN(n339), .Q(
        \bottom_add/A[10] ), .QN(n17) );
  DFFR_X1 \Data_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .RN(n339), .Q(
        \bottom_add/A[9] ), .QN(n18) );
  DFFR_X1 \dataBottom_reg[13]  ( .D(\U6/Z_13 ), .CK(clock), .RN(n339), .Q(
        \U4/DATA1_13 ) );
  DFFR_X1 \dataBottom_reg[12]  ( .D(\U6/Z_12 ), .CK(clock), .RN(n339), .Q(
        \U4/DATA1_12 ) );
  DFFR_X1 \dataBottom_reg[11]  ( .D(\U6/Z_11 ), .CK(clock), .RN(n339), .Q(
        \U4/DATA1_11 ) );
  DFFR_X1 \dataBottom_reg[10]  ( .D(\U6/Z_10 ), .CK(clock), .RN(n339), .Q(
        \U4/DATA1_10 ) );
  DFFR_X1 \dataBottom_reg[9]  ( .D(\U6/Z_9 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_9 ) );
  DFFR_X1 \dataBottom_reg[8]  ( .D(\U6/Z_8 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_8 ) );
  DFFR_X1 \dataBottom_reg[7]  ( .D(\U6/Z_7 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_7 ) );
  DFFR_X1 \dataBottom_reg[6]  ( .D(\U6/Z_6 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_6 ) );
  DFFR_X1 \dataBottom_reg[5]  ( .D(\U6/Z_5 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_5 ) );
  DFFR_X1 \dataBottom_reg[4]  ( .D(\U6/Z_4 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_4 ) );
  DFFR_X1 \dataBottom_reg[3]  ( .D(\U6/Z_3 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_3 ) );
  DFFR_X1 \dataBottom_reg[2]  ( .D(\U6/Z_2 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_2 ) );
  DFFR_X1 \dataBottom_reg[1]  ( .D(\U6/Z_1 ), .CK(clock), .RN(n340), .Q(
        \U4/DATA1_1 ) );
  DFFR_X1 dataCout_reg ( .D(\U5/Z_0 ), .CK(clock), .RN(n340), .Q(\top_add/CI ), 
        .QN(n312) );
  DFFR_X1 \dataTop_reg[18]  ( .D(\U8/Z_12 ), .CK(clock), .RN(n341), .Q(
        \top_add/A[12] ), .QN(n21) );
  DFFR_X1 \dataTop_reg[17]  ( .D(\U8/Z_11 ), .CK(clock), .RN(n341), .Q(
        \top_add/A[11] ), .QN(n22) );
  DFFR_X1 \dataTop_reg[16]  ( .D(\U8/Z_10 ), .CK(clock), .RN(n341), .Q(n309), 
        .QN(n23) );
  DFFR_X1 \dataTop_reg[15]  ( .D(\U8/Z_9 ), .CK(clock), .RN(n341), .Q(n305), 
        .QN(n24) );
  DFFR_X1 \dataTop_reg[14]  ( .D(\U8/Z_8 ), .CK(clock), .RN(n341), .Q(n306), 
        .QN(n25) );
  DFFR_X1 \DataOut_reg[27]  ( .D(\U4/Z_27 ), .CK(clock), .RN(n342), .Q(
        DataOut[27]) );
  DFFR_X1 \DataOut_reg[26]  ( .D(\U4/Z_26 ), .CK(clock), .RN(n342), .Q(
        DataOut[26]) );
  DFFR_X1 \DataOut_reg[25]  ( .D(\U4/Z_25 ), .CK(clock), .RN(n342), .Q(
        DataOut[25]) );
  DFFR_X1 \DataOut_reg[24]  ( .D(\U4/Z_24 ), .CK(clock), .RN(n342), .Q(
        DataOut[24]) );
  DFFR_X1 \DataOut_reg[23]  ( .D(\U4/Z_23 ), .CK(clock), .RN(n342), .Q(
        DataOut[23]) );
  DFFR_X1 \DataOut_reg[22]  ( .D(\U4/Z_22 ), .CK(clock), .RN(n342), .Q(
        DataOut[22]) );
  DFFR_X1 \DataOut_reg[21]  ( .D(\U4/Z_21 ), .CK(clock), .RN(n342), .Q(
        DataOut[21]) );
  DFFR_X1 \DataOut_reg[20]  ( .D(\U4/Z_20 ), .CK(clock), .RN(n342), .Q(
        DataOut[20]) );
  DFFR_X1 \DataOut_reg[19]  ( .D(\U4/Z_19 ), .CK(clock), .RN(n342), .Q(
        DataOut[19]) );
  DFFR_X1 \DataOut_reg[18]  ( .D(\U4/Z_18 ), .CK(clock), .RN(n343), .Q(
        DataOut[18]) );
  DFFR_X1 \DataOut_reg[17]  ( .D(\U4/Z_17 ), .CK(clock), .RN(n343), .Q(
        DataOut[17]) );
  DFFR_X1 \DataOut_reg[16]  ( .D(\U4/Z_16 ), .CK(clock), .RN(n343), .Q(
        DataOut[16]) );
  DFFR_X1 \DataOut_reg[15]  ( .D(\U4/Z_15 ), .CK(clock), .RN(n343), .Q(
        DataOut[15]) );
  DFFR_X1 \DataOut_reg[14]  ( .D(\U4/Z_14 ), .CK(clock), .RN(n343), .Q(
        DataOut[14]) );
  AND2_X1 U81 ( .A1(\U4/DATA1_6 ), .A2(n81), .ZN(\U4/Z_6 ) );
  AND2_X1 U82 ( .A1(\U4/DATA1_5 ), .A2(n81), .ZN(\U4/Z_5 ) );
  AND2_X1 U83 ( .A1(\U4/DATA1_4 ), .A2(n81), .ZN(\U4/Z_4 ) );
  AND2_X1 U84 ( .A1(\U4/DATA1_3 ), .A2(n81), .ZN(\U4/Z_3 ) );
  AND2_X1 U93 ( .A1(\U4/DATA1_2 ), .A2(n81), .ZN(\U4/Z_2 ) );
  AND2_X1 U104 ( .A1(\U4/DATA1_1 ), .A2(n81), .ZN(\U4/Z_1 ) );
  DFFR_X2 \Data_reg[19]  ( .D(\U7/Z_19 ), .CK(clock), .RN(reset_n), .Q(
        \U8/DATA1_13 ) );
  SDFFRS_X2 \Data_reg[0]  ( .D(1'b0), .SI(StartIn), .SE(\U7/DATA1_0 ), .CK(
        clock), .RN(n602), .SN(n603), .Q(\bottom_add/A[8] ), .QN(n311) );
  DFFR_X2 \dataBottom_reg[0]  ( .D(n316), .CK(clock), .RN(reset_n), .Q(
        \U4/DATA1_0 ) );
  DFFR_X2 \Data_reg[6]  ( .D(\U7/Z_6 ), .CK(clock), .RN(n339), .QN(n13) );
  DFFR_X2 \Data_reg[7]  ( .D(\U7/Z_7 ), .CK(clock), .RN(n339), .QN(n12) );
  DFFR_X2 \Data_reg[8]  ( .D(\U7/Z_8 ), .CK(clock), .RN(n339), .Q(n456), .QN(
        n11) );
  DFFR_X2 \Data_reg[9]  ( .D(\U7/Z_9 ), .CK(clock), .RN(n344), .Q(n465), .QN(
        n10) );
  DFFR_X2 \Data_reg[10]  ( .D(\U7/Z_10 ), .CK(clock), .RN(n340), .Q(n474), 
        .QN(n9) );
  DFFR_X2 \Data_reg[11]  ( .D(\U7/Z_11 ), .CK(clock), .RN(n344), .Q(n483), 
        .QN(n8) );
  DFFR_X2 \Data_reg[12]  ( .D(\U7/Z_12 ), .CK(clock), .RN(n340), .Q(n492), 
        .QN(n7) );
  DFFR_X2 \Data_reg[13]  ( .D(\U7/Z_13 ), .CK(clock), .RN(n344), .Q(n498), 
        .QN(n6) );
  DFFR_X2 Start0_reg ( .D(StartIn), .CK(clock), .RN(reset_n), .Q(n162), .QN(
        n600) );
  DFFR_X2 \dataTop_reg[19]  ( .D(\U8/Z_13 ), .CK(clock), .RN(reset_n), .Q(
        \top_add/A[13] ), .QN(n20) );
  DFFR_X2 \dataTop_reg[7]  ( .D(\U8/Z_1 ), .CK(clock), .RN(n342), .Q(
        \top_add/A[1] ), .QN(n517) );
  DFFR_X2 \dataTop_reg[6]  ( .D(\U8/Z_0 ), .CK(clock), .RN(n342), .Q(
        \top_add/A[0] ), .QN(n508) );
  DFFR_X2 \dataTop_reg[8]  ( .D(\U8/Z_2 ), .CK(clock), .RN(n341), .Q(
        \top_add/A[2] ), .QN(n527) );
  DFFR_X2 \dataTop_reg[13]  ( .D(\U8/Z_7 ), .CK(clock), .RN(n341), .QN(n571)
         );
  DFFR_X2 \dataTop_reg[12]  ( .D(\U8/Z_6 ), .CK(clock), .RN(n341), .QN(n567)
         );
  DFFR_X2 \dataTop_reg[11]  ( .D(\U8/Z_5 ), .CK(clock), .RN(n341), .Q(
        \top_add/A[5] ), .QN(n565) );
  DFFR_X2 \dataTop_reg[10]  ( .D(\U8/Z_4 ), .CK(clock), .RN(n341), .Q(
        \top_add/A[4] ), .QN(n559) );
  DFFR_X2 \dataTop_reg[9]  ( .D(\U8/Z_3 ), .CK(clock), .RN(n341), .Q(
        \top_add/A[3] ), .QN(n545) );
  DFFR_X2 \DataOut_reg[13]  ( .D(\U4/Z_13 ), .CK(clock), .RN(n343), .Q(
        DataOut[13]) );
  DFFR_X2 \DataOut_reg[12]  ( .D(\U4/Z_12 ), .CK(clock), .RN(n343), .Q(
        DataOut[12]) );
  DFFR_X2 \DataOut_reg[11]  ( .D(\U4/Z_11 ), .CK(clock), .RN(n343), .Q(
        DataOut[11]) );
  DFFR_X2 \DataOut_reg[10]  ( .D(\U4/Z_10 ), .CK(clock), .RN(n343), .Q(
        DataOut[10]) );
  DFFR_X2 \DataOut_reg[9]  ( .D(\U4/Z_9 ), .CK(clock), .RN(n343), .Q(
        DataOut[9]) );
  DFFR_X2 \DataOut_reg[8]  ( .D(\U4/Z_8 ), .CK(clock), .RN(n343), .Q(
        DataOut[8]) );
  DFFR_X2 \DataOut_reg[7]  ( .D(\U4/Z_7 ), .CK(clock), .RN(n343), .Q(
        DataOut[7]) );
  DFFR_X2 \DataOut_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n344), .Q(
        DataOut[6]) );
  DFFR_X2 \DataOut_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n344), .Q(
        DataOut[5]) );
  DFFR_X2 \DataOut_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(n344), .Q(
        DataOut[4]) );
  DFFR_X2 \DataOut_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n344), .Q(
        DataOut[3]) );
  DFFR_X2 \DataOut_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .RN(n344), .Q(
        DataOut[2]) );
  DFFR_X2 \DataOut_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .RN(n344), .Q(
        DataOut[1]) );
  DFFR_X2 \DataOut_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n340), .Q(
        DataOut[0]) );
  DFFR_X2 Start1_reg ( .D(n162), .CK(clock), .RN(reset_n), .Q(n81), .QN(n587)
         );
  DFFR_X2 StartOut_reg ( .D(n81), .CK(clock), .RN(n342), .Q(StartOut) );
  DFFR_X2 \Data_reg[14]  ( .D(\U7/Z_14 ), .CK(clock), .RN(n344), .Q(
        \U8/DATA1_8 ) );
  DFFR_X2 \Data_reg[16]  ( .D(\U7/Z_16 ), .CK(clock), .RN(n340), .Q(
        \U8/DATA1_10 ) );
  DFFR_X2 \Data_reg[18]  ( .D(\U7/Z_18 ), .CK(clock), .RN(n344), .Q(
        \U8/DATA1_12 ) );
  DFFR_X2 \Data_reg[15]  ( .D(\U7/Z_15 ), .CK(clock), .RN(n344), .Q(
        \U8/DATA1_9 ) );
  DFFR_X2 \Data_reg[17]  ( .D(\U7/Z_17 ), .CK(clock), .RN(n344), .Q(
        \U8/DATA1_11 ) );
  OAI221_X2 U3 ( .B1(n555), .B2(n338), .C1(n556), .C2(n552), .A(n337), .ZN(
        n336) );
  INV_X1 U4 ( .A(n556), .ZN(n555) );
  AOI211_X2 U5 ( .C1(n399), .C2(n398), .A(n397), .B(n396), .ZN(n407) );
  AOI22_X2 U7 ( .A1(n433), .A2(n432), .B1(\first_add/A[15] ), .B2(n431), .ZN(
        n513) );
  NOR2_X2 U8 ( .A1(\first_add/A[1] ), .A2(n347), .ZN(n348) );
  INV_X4 U9 ( .A(n487), .ZN(n426) );
  BUF_X4 U10 ( .A(n377), .Z(n327) );
  AND2_X4 U11 ( .A1(n308), .A2(n25), .ZN(n304) );
  AND2_X4 U12 ( .A1(n304), .A2(n24), .ZN(n307) );
  AND2_X4 U13 ( .A1(n313), .A2(n571), .ZN(n308) );
  XNOR2_X2 U14 ( .A(n531), .B(CdfMin[18]), .ZN(n310) );
  AND2_X4 U15 ( .A1(n568), .A2(n567), .ZN(n313) );
  AND2_X4 U16 ( .A1(n402), .A2(n400), .ZN(n314) );
  XNOR2_X2 U17 ( .A(n549), .B(CdfMin[19]), .ZN(n315) );
  AND2_X1 U18 ( .A1(\bottom_add/A[8] ), .A2(n162), .ZN(n316) );
  NAND2_X1 U19 ( .A1(n537), .A2(n522), .ZN(n317) );
  XNOR2_X2 U20 ( .A(n318), .B(n326), .ZN(n514) );
  XOR2_X2 U21 ( .A(CdfMin[16]), .B(\first_add/A[16] ), .Z(n318) );
  NAND2_X2 U22 ( .A1(n401), .A2(n314), .ZN(n406) );
  NAND2_X2 U23 ( .A1(n351), .A2(n375), .ZN(n323) );
  NAND2_X1 U24 ( .A1(\first_add/A[3] ), .A2(n353), .ZN(n393) );
  NAND2_X1 U25 ( .A1(n354), .A2(n393), .ZN(n357) );
  INV_X1 U26 ( .A(n353), .ZN(n319) );
  AND2_X4 U27 ( .A1(n400), .A2(n402), .ZN(n399) );
  NAND2_X2 U28 ( .A1(CdfMin[4]), .A2(n356), .ZN(n400) );
  NOR2_X2 U29 ( .A1(n320), .A2(\first_add/A[0] ), .ZN(n322) );
  INV_X4 U30 ( .A(CdfMin[0]), .ZN(n320) );
  INV_X1 U31 ( .A(n460), .ZN(n461) );
  INV_X1 U32 ( .A(n322), .ZN(n383) );
  OR2_X4 U33 ( .A1(n353), .A2(\first_add/A[3] ), .ZN(n351) );
  NAND2_X1 U34 ( .A1(\first_add/A[0] ), .A2(n320), .ZN(n382) );
  INV_X8 U35 ( .A(n453), .ZN(n414) );
  AOI22_X2 U36 ( .A1(n417), .A2(n418), .B1(\first_add/A[10] ), .B2(n416), .ZN(
        n469) );
  INV_X1 U37 ( .A(n352), .ZN(n321) );
  INV_X1 U38 ( .A(CdfMin[4]), .ZN(n352) );
  XOR2_X1 U39 ( .A(n380), .B(n322), .Z(n381) );
  NAND3_X1 U40 ( .A1(n357), .A2(n402), .A3(n400), .ZN(n359) );
  NAND2_X1 U41 ( .A1(n372), .A2(n400), .ZN(n369) );
  NAND2_X1 U42 ( .A1(n383), .A2(n382), .ZN(\U7/DATA1_0 ) );
  INV_X2 U43 ( .A(CdfMin[6]), .ZN(n361) );
  NAND2_X1 U44 ( .A1(CdfMin[6]), .A2(n360), .ZN(n403) );
  INV_X1 U45 ( .A(CdfMin[5]), .ZN(n358) );
  NAND2_X1 U46 ( .A1(n359), .A2(n395), .ZN(n365) );
  INV_X2 U47 ( .A(n395), .ZN(n396) );
  OAI22_X2 U48 ( .A1(CdfMin[1]), .A2(n379), .B1(n322), .B2(n348), .ZN(n377) );
  NAND2_X2 U49 ( .A1(n324), .A2(CdfMin[2]), .ZN(n325) );
  NAND2_X2 U50 ( .A1(n325), .A2(n377), .ZN(n349) );
  INV_X4 U51 ( .A(\first_add/A[2] ), .ZN(n324) );
  XNOR2_X1 U52 ( .A(CdfMin[6]), .B(\first_add/A[6] ), .ZN(n366) );
  INV_X4 U53 ( .A(n394), .ZN(n397) );
  NAND2_X1 U54 ( .A1(n362), .A2(n394), .ZN(n363) );
  INV_X1 U55 ( .A(n505), .ZN(n506) );
  INV_X1 U56 ( .A(n500), .ZN(n501) );
  INV_X1 U57 ( .A(n478), .ZN(n479) );
  INV_X1 U58 ( .A(n487), .ZN(n488) );
  AOI22_X1 U59 ( .A1(n433), .A2(n432), .B1(\first_add/A[15] ), .B2(n431), .ZN(
        n326) );
  INV_X1 U60 ( .A(n420), .ZN(n328) );
  INV_X1 U61 ( .A(n446), .ZN(n447) );
  XNOR2_X1 U62 ( .A(n374), .B(n319), .ZN(n331) );
  XOR2_X1 U63 ( .A(n331), .B(n375), .Z(n376) );
  XOR2_X1 U64 ( .A(n329), .B(n327), .Z(n378) );
  XNOR2_X1 U65 ( .A(n324), .B(CdfMin[2]), .ZN(n329) );
  INV_X1 U66 ( .A(CdfMin[2]), .ZN(n346) );
  AND2_X2 U67 ( .A1(\first_add/A[7] ), .A2(n408), .ZN(n332) );
  AOI22_X4 U68 ( .A1(n421), .A2(n420), .B1(\first_add/A[11] ), .B2(n419), .ZN(
        n478) );
  AOI22_X4 U69 ( .A1(n424), .A2(n423), .B1(\first_add/A[12] ), .B2(n422), .ZN(
        n487) );
  AOI22_X4 U70 ( .A1(n426), .A2(n427), .B1(\first_add/A[13] ), .B2(n425), .ZN(
        n500) );
  AOI22_X4 U71 ( .A1(n429), .A2(n430), .B1(\first_add/A[14] ), .B2(n428), .ZN(
        n505) );
  AOI22_X4 U72 ( .A1(n414), .A2(n415), .B1(\first_add/A[9] ), .B2(n413), .ZN(
        n460) );
  XOR2_X1 U73 ( .A(\first_add/A[4] ), .B(n321), .Z(n335) );
  XNOR2_X1 U74 ( .A(CdfMin[7]), .B(\first_add/A[7] ), .ZN(n334) );
  XNOR2_X1 U75 ( .A(CdfMin[5]), .B(\first_add/A[5] ), .ZN(n333) );
  AOI211_X2 U76 ( .C1(n406), .C2(n407), .A(n405), .B(n404), .ZN(n409) );
  INV_X4 U77 ( .A(n345), .ZN(n344) );
  INV_X4 U78 ( .A(n345), .ZN(n341) );
  INV_X4 U79 ( .A(n345), .ZN(n340) );
  INV_X4 U80 ( .A(n345), .ZN(n343) );
  INV_X4 U85 ( .A(n345), .ZN(n342) );
  INV_X4 U86 ( .A(n345), .ZN(n339) );
  INV_X4 U87 ( .A(reset_n), .ZN(n345) );
  NAND2_X2 U88 ( .A1(n323), .A2(n368), .ZN(n401) );
  XNOR2_X2 U89 ( .A(n330), .B(n535), .ZN(n524) );
  XNOR2_X2 U90 ( .A(n521), .B(CdfMin[17]), .ZN(n330) );
  INV_X4 U91 ( .A(n336), .ZN(\U7/Z_19 ) );
  INV_X4 U92 ( .A(n554), .ZN(n337) );
  AND2_X1 U94 ( .A1(n435), .A2(CdfMin[16]), .ZN(n434) );
  AOI21_X2 U95 ( .B1(n584), .B2(n582), .A(n587), .ZN(\U4/Z_25 ) );
  XNOR2_X2 U96 ( .A(n370), .B(n333), .ZN(n371) );
  XNOR2_X2 U97 ( .A(n363), .B(n334), .ZN(n364) );
  XOR2_X2 U98 ( .A(n335), .B(n372), .Z(n373) );
  INV_X4 U99 ( .A(StartIn), .ZN(n523) );
  OR2_X4 U100 ( .A1(n550), .A2(n315), .ZN(n338) );
  INV_X1 U101 ( .A(n401), .ZN(n354) );
  NAND2_X1 U102 ( .A1(n323), .A2(n393), .ZN(n372) );
  NOR2_X1 U103 ( .A1(n310), .A2(n317), .ZN(n533) );
  NAND2_X1 U105 ( .A1(n551), .A2(n556), .ZN(n437) );
  INV_X2 U106 ( .A(n328), .ZN(n470) );
  INV_X2 U107 ( .A(n522), .ZN(n535) );
  NOR2_X4 U108 ( .A1(n409), .A2(n332), .ZN(n446) );
  INV_X4 U109 ( .A(\first_add/A[3] ), .ZN(n374) );
  NAND2_X2 U110 ( .A1(\first_add/A[2] ), .A2(n346), .ZN(n350) );
  INV_X4 U111 ( .A(\first_add/A[1] ), .ZN(n379) );
  INV_X4 U112 ( .A(CdfMin[1]), .ZN(n347) );
  NAND2_X2 U113 ( .A1(n350), .A2(n349), .ZN(n375) );
  NAND2_X2 U114 ( .A1(\first_add/A[4] ), .A2(n352), .ZN(n368) );
  INV_X4 U115 ( .A(CdfMin[3]), .ZN(n353) );
  INV_X4 U116 ( .A(\first_add/A[5] ), .ZN(n355) );
  NAND2_X2 U117 ( .A1(CdfMin[5]), .A2(n355), .ZN(n402) );
  INV_X4 U118 ( .A(\first_add/A[4] ), .ZN(n356) );
  NAND2_X2 U119 ( .A1(\first_add/A[5] ), .A2(n358), .ZN(n395) );
  INV_X4 U120 ( .A(\first_add/A[6] ), .ZN(n360) );
  NAND2_X2 U121 ( .A1(n365), .A2(n403), .ZN(n362) );
  NAND2_X2 U122 ( .A1(n361), .A2(\first_add/A[6] ), .ZN(n394) );
  NOR2_X2 U123 ( .A1(n364), .A2(n523), .ZN(\U7/Z_7 ) );
  XNOR2_X2 U124 ( .A(n366), .B(n365), .ZN(n367) );
  NOR2_X2 U125 ( .A1(n367), .A2(n523), .ZN(\U7/Z_6 ) );
  NAND2_X2 U126 ( .A1(n369), .A2(n368), .ZN(n370) );
  NOR2_X2 U127 ( .A1(n371), .A2(n523), .ZN(\U7/Z_5 ) );
  NOR2_X2 U128 ( .A1(n373), .A2(n523), .ZN(\U7/Z_4 ) );
  NOR2_X2 U129 ( .A1(n376), .A2(n523), .ZN(\U7/Z_3 ) );
  NOR2_X2 U130 ( .A1(n378), .A2(n523), .ZN(\U7/Z_2 ) );
  XOR2_X2 U131 ( .A(n379), .B(CdfMin[1]), .Z(n380) );
  NOR2_X2 U132 ( .A1(n381), .A2(n523), .ZN(\U7/Z_1 ) );
  INV_X4 U133 ( .A(\first_add/A[18] ), .ZN(n531) );
  NAND2_X2 U134 ( .A1(CdfMin[18]), .A2(n531), .ZN(n551) );
  INV_X4 U135 ( .A(CdfMin[17]), .ZN(n384) );
  NAND2_X2 U136 ( .A1(\first_add/A[17] ), .A2(n384), .ZN(n536) );
  INV_X4 U137 ( .A(\first_add/A[17] ), .ZN(n521) );
  NAND2_X2 U138 ( .A1(CdfMin[17]), .A2(n521), .ZN(n537) );
  INV_X4 U139 ( .A(\first_add/A[16] ), .ZN(n435) );
  INV_X4 U140 ( .A(\first_add/A[15] ), .ZN(n385) );
  NAND2_X2 U141 ( .A1(CdfMin[15]), .A2(n385), .ZN(n433) );
  INV_X4 U142 ( .A(\first_add/A[14] ), .ZN(n386) );
  NAND2_X2 U143 ( .A1(CdfMin[14]), .A2(n386), .ZN(n430) );
  INV_X4 U144 ( .A(\first_add/A[13] ), .ZN(n387) );
  NAND2_X2 U145 ( .A1(CdfMin[13]), .A2(n387), .ZN(n427) );
  INV_X4 U146 ( .A(\first_add/A[12] ), .ZN(n388) );
  NAND2_X2 U147 ( .A1(CdfMin[12]), .A2(n388), .ZN(n424) );
  INV_X4 U148 ( .A(\first_add/A[11] ), .ZN(n389) );
  NAND2_X2 U149 ( .A1(CdfMin[11]), .A2(n389), .ZN(n421) );
  INV_X4 U150 ( .A(\first_add/A[10] ), .ZN(n390) );
  NAND2_X2 U151 ( .A1(CdfMin[10]), .A2(n390), .ZN(n418) );
  INV_X4 U152 ( .A(\first_add/A[9] ), .ZN(n391) );
  NAND2_X2 U153 ( .A1(CdfMin[9]), .A2(n391), .ZN(n415) );
  INV_X4 U154 ( .A(\first_add/A[8] ), .ZN(n392) );
  NAND2_X2 U155 ( .A1(CdfMin[8]), .A2(n392), .ZN(n412) );
  INV_X4 U156 ( .A(n393), .ZN(n398) );
  INV_X4 U157 ( .A(n403), .ZN(n405) );
  INV_X4 U158 ( .A(CdfMin[7]), .ZN(n408) );
  NOR2_X2 U159 ( .A1(\first_add/A[7] ), .A2(n408), .ZN(n404) );
  INV_X4 U160 ( .A(n446), .ZN(n411) );
  INV_X4 U161 ( .A(CdfMin[8]), .ZN(n410) );
  AOI22_X4 U162 ( .A1(n411), .A2(n412), .B1(\first_add/A[8] ), .B2(n410), .ZN(
        n453) );
  INV_X4 U163 ( .A(CdfMin[9]), .ZN(n413) );
  INV_X4 U164 ( .A(n460), .ZN(n417) );
  INV_X4 U165 ( .A(CdfMin[10]), .ZN(n416) );
  INV_X4 U166 ( .A(n469), .ZN(n420) );
  INV_X4 U167 ( .A(CdfMin[11]), .ZN(n419) );
  INV_X4 U168 ( .A(n478), .ZN(n423) );
  INV_X4 U169 ( .A(CdfMin[12]), .ZN(n422) );
  INV_X4 U170 ( .A(CdfMin[13]), .ZN(n425) );
  INV_X4 U171 ( .A(n500), .ZN(n429) );
  INV_X4 U172 ( .A(CdfMin[14]), .ZN(n428) );
  INV_X4 U173 ( .A(n505), .ZN(n432) );
  INV_X4 U174 ( .A(CdfMin[15]), .ZN(n431) );
  OAI22_X2 U175 ( .A1(CdfMin[16]), .A2(n435), .B1(n513), .B2(n434), .ZN(n522)
         );
  NAND2_X2 U176 ( .A1(n522), .A2(n537), .ZN(n532) );
  NAND2_X2 U177 ( .A1(n532), .A2(n536), .ZN(n556) );
  INV_X4 U178 ( .A(CdfMin[18]), .ZN(n436) );
  NAND2_X2 U179 ( .A1(\first_add/A[18] ), .A2(n436), .ZN(n553) );
  NAND2_X2 U180 ( .A1(n437), .A2(n553), .ZN(n440) );
  INV_X4 U181 ( .A(\first_add/A[19] ), .ZN(n549) );
  NAND2_X2 U182 ( .A1(CdfMin[19]), .A2(n549), .ZN(n443) );
  NAND2_X2 U183 ( .A1(n440), .A2(n443), .ZN(n439) );
  INV_X4 U184 ( .A(CdfMin[19]), .ZN(n438) );
  NAND2_X2 U185 ( .A1(\first_add/A[19] ), .A2(n438), .ZN(n441) );
  NAND3_X2 U186 ( .A1(n439), .A2(n345), .A3(n441), .ZN(n602) );
  INV_X4 U187 ( .A(n440), .ZN(n442) );
  NAND2_X2 U188 ( .A1(n442), .A2(n441), .ZN(n444) );
  NAND3_X2 U189 ( .A1(n444), .A2(n443), .A3(n345), .ZN(n603) );
  NAND3_X2 U190 ( .A1(n18), .A2(n17), .A3(n311), .ZN(n591) );
  INV_X4 U191 ( .A(n591), .ZN(n593) );
  NAND3_X2 U192 ( .A1(n16), .A2(n15), .A3(n593), .ZN(n596) );
  INV_X4 U193 ( .A(n596), .ZN(n598) );
  NAND3_X2 U194 ( .A1(n13), .A2(n14), .A3(n598), .ZN(n449) );
  XOR2_X2 U195 ( .A(n449), .B(n12), .Z(n445) );
  NOR2_X2 U196 ( .A1(n600), .A2(n445), .ZN(\U6/Z_7 ) );
  AND2_X1 U197 ( .A1(\U4/DATA1_7 ), .A2(n81), .ZN(\U4/Z_7 ) );
  FA_X1 U198 ( .A(\first_add/A[8] ), .B(CdfMin[8]), .CI(n447), .S(n448) );
  NOR2_X2 U199 ( .A1(n448), .A2(n523), .ZN(\U7/Z_8 ) );
  XNOR2_X2 U200 ( .A(n11), .B(\bottom_add/A[8] ), .ZN(n451) );
  INV_X4 U201 ( .A(n449), .ZN(n450) );
  NAND2_X2 U202 ( .A1(n12), .A2(n450), .ZN(n455) );
  XNOR2_X2 U203 ( .A(n451), .B(n455), .ZN(n452) );
  NOR2_X2 U204 ( .A1(n452), .A2(n600), .ZN(\U6/Z_8 ) );
  AND2_X1 U205 ( .A1(\U4/DATA1_8 ), .A2(n81), .ZN(\U4/Z_8 ) );
  FA_X1 U206 ( .A(\first_add/A[9] ), .B(CdfMin[9]), .CI(n414), .S(n454) );
  NOR2_X2 U207 ( .A1(n454), .A2(n523), .ZN(\U7/Z_9 ) );
  OAI22_X2 U208 ( .A1(n456), .A2(n311), .B1(n455), .B2(n456), .ZN(n457) );
  INV_X4 U209 ( .A(n457), .ZN(n464) );
  XOR2_X2 U210 ( .A(\bottom_add/A[9] ), .B(n10), .Z(n458) );
  XOR2_X2 U211 ( .A(n464), .B(n458), .Z(n459) );
  NOR2_X2 U212 ( .A1(n459), .A2(n600), .ZN(\U6/Z_9 ) );
  AND2_X1 U213 ( .A1(\U4/DATA1_9 ), .A2(n81), .ZN(\U4/Z_9 ) );
  FA_X1 U214 ( .A(\first_add/A[10] ), .B(CdfMin[10]), .CI(n461), .S(n462) );
  NOR2_X2 U215 ( .A1(n462), .A2(n523), .ZN(\U7/Z_10 ) );
  NOR2_X2 U216 ( .A1(\bottom_add/A[9] ), .A2(n10), .ZN(n463) );
  OAI22_X2 U217 ( .A1(n465), .A2(n18), .B1(n464), .B2(n463), .ZN(n466) );
  INV_X4 U218 ( .A(n466), .ZN(n473) );
  XOR2_X2 U219 ( .A(\bottom_add/A[10] ), .B(n9), .Z(n467) );
  XOR2_X2 U220 ( .A(n473), .B(n467), .Z(n468) );
  NOR2_X2 U221 ( .A1(n468), .A2(n600), .ZN(\U6/Z_10 ) );
  AND2_X1 U222 ( .A1(\U4/DATA1_10 ), .A2(n81), .ZN(\U4/Z_10 ) );
  FA_X1 U223 ( .A(\first_add/A[11] ), .B(CdfMin[11]), .CI(n470), .S(n471) );
  NOR2_X2 U224 ( .A1(n471), .A2(n523), .ZN(\U7/Z_11 ) );
  NOR2_X2 U225 ( .A1(\bottom_add/A[10] ), .A2(n9), .ZN(n472) );
  OAI22_X2 U226 ( .A1(n474), .A2(n17), .B1(n473), .B2(n472), .ZN(n475) );
  INV_X4 U227 ( .A(n475), .ZN(n482) );
  XOR2_X2 U228 ( .A(\bottom_add/A[11] ), .B(n8), .Z(n476) );
  XOR2_X2 U229 ( .A(n482), .B(n476), .Z(n477) );
  NOR2_X2 U230 ( .A1(n477), .A2(n600), .ZN(\U6/Z_11 ) );
  AND2_X1 U231 ( .A1(\U4/DATA1_11 ), .A2(n81), .ZN(\U4/Z_11 ) );
  FA_X1 U232 ( .A(\first_add/A[12] ), .B(CdfMin[12]), .CI(n479), .S(n480) );
  NOR2_X2 U233 ( .A1(n480), .A2(n523), .ZN(\U7/Z_12 ) );
  NOR2_X2 U234 ( .A1(\bottom_add/A[11] ), .A2(n8), .ZN(n481) );
  OAI22_X2 U235 ( .A1(n483), .A2(n16), .B1(n482), .B2(n481), .ZN(n484) );
  INV_X4 U236 ( .A(n484), .ZN(n491) );
  XOR2_X2 U237 ( .A(\bottom_add/A[12] ), .B(n7), .Z(n485) );
  XOR2_X2 U238 ( .A(n491), .B(n485), .Z(n486) );
  NOR2_X2 U239 ( .A1(n486), .A2(n600), .ZN(\U6/Z_12 ) );
  AND2_X1 U240 ( .A1(\U4/DATA1_12 ), .A2(n81), .ZN(\U4/Z_12 ) );
  FA_X1 U241 ( .A(\first_add/A[13] ), .B(CdfMin[13]), .CI(n488), .S(n489) );
  NOR2_X2 U242 ( .A1(n489), .A2(n523), .ZN(\U7/Z_13 ) );
  NOR2_X2 U243 ( .A1(\bottom_add/A[12] ), .A2(n7), .ZN(n490) );
  OAI22_X2 U244 ( .A1(n492), .A2(n15), .B1(n491), .B2(n490), .ZN(n493) );
  INV_X4 U245 ( .A(n493), .ZN(n497) );
  XOR2_X2 U246 ( .A(\bottom_add/A[13] ), .B(n6), .Z(n494) );
  XOR2_X2 U247 ( .A(n497), .B(n494), .Z(n495) );
  NOR2_X2 U248 ( .A1(n495), .A2(n600), .ZN(\U6/Z_13 ) );
  AND2_X1 U249 ( .A1(\U4/DATA1_13 ), .A2(n81), .ZN(\U4/Z_13 ) );
  NOR2_X2 U250 ( .A1(\bottom_add/A[13] ), .A2(n6), .ZN(n496) );
  OAI22_X2 U251 ( .A1(n498), .A2(n14), .B1(n497), .B2(n496), .ZN(n499) );
  AND2_X1 U252 ( .A1(n162), .A2(n499), .ZN(\U5/Z_0 ) );
  FA_X1 U253 ( .A(\first_add/A[14] ), .B(CdfMin[14]), .CI(n501), .S(n502) );
  NOR2_X2 U254 ( .A1(n502), .A2(n523), .ZN(\U7/Z_14 ) );
  AND2_X1 U255 ( .A1(\U8/DATA1_8 ), .A2(n162), .ZN(\U8/Z_8 ) );
  NOR2_X2 U256 ( .A1(n600), .A2(n13), .ZN(\U8/Z_0 ) );
  XOR2_X2 U257 ( .A(n312), .B(n25), .Z(n503) );
  XOR2_X2 U258 ( .A(n503), .B(\top_add/A[0] ), .Z(n504) );
  NOR2_X2 U259 ( .A1(n504), .A2(n587), .ZN(\U4/Z_14 ) );
  FA_X1 U260 ( .A(\first_add/A[15] ), .B(CdfMin[15]), .CI(n506), .S(n507) );
  NOR2_X2 U261 ( .A1(n507), .A2(n523), .ZN(\U7/Z_15 ) );
  AND2_X1 U262 ( .A1(\U8/DATA1_9 ), .A2(n162), .ZN(\U8/Z_9 ) );
  NOR2_X2 U263 ( .A1(n600), .A2(n12), .ZN(\U8/Z_1 ) );
  NOR2_X2 U264 ( .A1(n25), .A2(\top_add/CI ), .ZN(n509) );
  OAI22_X2 U265 ( .A1(n312), .A2(n306), .B1(n509), .B2(n508), .ZN(n510) );
  INV_X4 U266 ( .A(n510), .ZN(n516) );
  XOR2_X2 U267 ( .A(\top_add/A[1] ), .B(n24), .Z(n511) );
  XOR2_X2 U268 ( .A(n516), .B(n511), .Z(n512) );
  NOR2_X2 U269 ( .A1(n512), .A2(n587), .ZN(\U4/Z_15 ) );
  NOR2_X2 U270 ( .A1(n514), .A2(n523), .ZN(\U7/Z_16 ) );
  AND2_X1 U271 ( .A1(\U8/DATA1_10 ), .A2(n162), .ZN(\U8/Z_10 ) );
  NOR2_X2 U272 ( .A1(n600), .A2(n11), .ZN(\U8/Z_2 ) );
  NOR2_X2 U273 ( .A1(\top_add/A[1] ), .A2(n24), .ZN(n515) );
  OAI22_X2 U274 ( .A1(n305), .A2(n517), .B1(n516), .B2(n515), .ZN(n518) );
  INV_X4 U275 ( .A(n518), .ZN(n526) );
  XOR2_X2 U276 ( .A(\top_add/A[2] ), .B(n23), .Z(n519) );
  XOR2_X2 U277 ( .A(n526), .B(n519), .Z(n520) );
  NOR2_X2 U278 ( .A1(n520), .A2(n587), .ZN(\U4/Z_16 ) );
  NOR2_X2 U279 ( .A1(n524), .A2(n523), .ZN(\U7/Z_17 ) );
  AND2_X1 U280 ( .A1(\U8/DATA1_11 ), .A2(n162), .ZN(\U8/Z_11 ) );
  NOR2_X2 U281 ( .A1(n600), .A2(n10), .ZN(\U8/Z_3 ) );
  NOR2_X2 U282 ( .A1(\top_add/A[2] ), .A2(n23), .ZN(n525) );
  OAI22_X2 U283 ( .A1(n309), .A2(n527), .B1(n526), .B2(n525), .ZN(n528) );
  INV_X4 U284 ( .A(n528), .ZN(n544) );
  XOR2_X2 U285 ( .A(\top_add/A[3] ), .B(n22), .Z(n529) );
  XOR2_X2 U286 ( .A(n544), .B(n529), .Z(n530) );
  NOR2_X2 U287 ( .A1(n530), .A2(n587), .ZN(\U4/Z_17 ) );
  NOR2_X2 U288 ( .A1(n310), .A2(n536), .ZN(n534) );
  NOR2_X2 U289 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND3_X2 U290 ( .A1(n536), .A2(n310), .A3(n535), .ZN(n540) );
  INV_X4 U291 ( .A(n537), .ZN(n538) );
  NAND2_X2 U292 ( .A1(n538), .A2(n310), .ZN(n539) );
  NAND4_X2 U293 ( .A1(n541), .A2(n540), .A3(n539), .A4(StartIn), .ZN(n542) );
  INV_X4 U294 ( .A(n542), .ZN(\U7/Z_18 ) );
  AND2_X1 U295 ( .A1(\U8/DATA1_12 ), .A2(n162), .ZN(\U8/Z_12 ) );
  NOR2_X2 U296 ( .A1(n600), .A2(n9), .ZN(\U8/Z_4 ) );
  NOR2_X2 U297 ( .A1(\top_add/A[3] ), .A2(n22), .ZN(n543) );
  OAI22_X2 U298 ( .A1(\top_add/A[11] ), .A2(n545), .B1(n544), .B2(n543), .ZN(
        n546) );
  INV_X4 U299 ( .A(n546), .ZN(n558) );
  XOR2_X2 U300 ( .A(\top_add/A[4] ), .B(n21), .Z(n547) );
  XOR2_X2 U301 ( .A(n558), .B(n547), .Z(n548) );
  NOR2_X2 U302 ( .A1(n548), .A2(n587), .ZN(\U4/Z_18 ) );
  INV_X4 U303 ( .A(n551), .ZN(n550) );
  NAND2_X2 U304 ( .A1(n553), .A2(n315), .ZN(n552) );
  OAI221_X2 U305 ( .B1(n315), .B2(n553), .C1(n552), .C2(n551), .A(StartIn), 
        .ZN(n554) );
  AND2_X1 U306 ( .A1(\U8/DATA1_13 ), .A2(n162), .ZN(\U8/Z_13 ) );
  NOR2_X2 U307 ( .A1(n600), .A2(n8), .ZN(\U8/Z_5 ) );
  NOR2_X2 U308 ( .A1(\top_add/A[4] ), .A2(n21), .ZN(n557) );
  OAI22_X2 U309 ( .A1(\top_add/A[12] ), .A2(n559), .B1(n558), .B2(n557), .ZN(
        n560) );
  INV_X4 U310 ( .A(n560), .ZN(n564) );
  XOR2_X2 U311 ( .A(\top_add/A[5] ), .B(n20), .Z(n561) );
  XOR2_X2 U312 ( .A(n564), .B(n561), .Z(n562) );
  NOR2_X2 U313 ( .A1(n562), .A2(n587), .ZN(\U4/Z_19 ) );
  NOR2_X2 U314 ( .A1(n600), .A2(n7), .ZN(\U8/Z_6 ) );
  NOR2_X2 U315 ( .A1(\top_add/A[5] ), .A2(n20), .ZN(n563) );
  OAI22_X2 U316 ( .A1(\top_add/A[13] ), .A2(n565), .B1(n564), .B2(n563), .ZN(
        n566) );
  INV_X4 U317 ( .A(n566), .ZN(n568) );
  NOR2_X2 U318 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X2 U319 ( .A1(n313), .A2(n569), .ZN(n570) );
  NOR2_X2 U320 ( .A1(n570), .A2(n587), .ZN(\U4/Z_20 ) );
  NOR2_X2 U321 ( .A1(n600), .A2(n6), .ZN(\U8/Z_7 ) );
  NOR2_X2 U322 ( .A1(n313), .A2(n571), .ZN(n572) );
  NOR2_X2 U323 ( .A1(n308), .A2(n572), .ZN(n573) );
  NOR2_X2 U324 ( .A1(n573), .A2(n587), .ZN(\U4/Z_21 ) );
  NOR2_X2 U325 ( .A1(n308), .A2(n25), .ZN(n574) );
  NOR2_X2 U326 ( .A1(n304), .A2(n574), .ZN(n575) );
  NOR2_X2 U327 ( .A1(n575), .A2(n587), .ZN(\U4/Z_22 ) );
  NOR2_X2 U328 ( .A1(n304), .A2(n24), .ZN(n576) );
  NOR2_X2 U329 ( .A1(n307), .A2(n576), .ZN(n577) );
  NOR2_X2 U330 ( .A1(n577), .A2(n587), .ZN(\U4/Z_23 ) );
  NAND2_X2 U331 ( .A1(n307), .A2(n23), .ZN(n581) );
  INV_X4 U332 ( .A(n581), .ZN(n580) );
  NOR2_X2 U333 ( .A1(n307), .A2(n23), .ZN(n578) );
  NOR2_X2 U334 ( .A1(n580), .A2(n578), .ZN(n579) );
  NOR2_X2 U335 ( .A1(n579), .A2(n587), .ZN(\U4/Z_24 ) );
  NAND2_X2 U336 ( .A1(n580), .A2(n22), .ZN(n584) );
  NAND2_X2 U337 ( .A1(\top_add/A[11] ), .A2(n581), .ZN(n582) );
  XOR2_X2 U338 ( .A(n584), .B(\top_add/A[12] ), .Z(n583) );
  NOR2_X2 U339 ( .A1(n587), .A2(n583), .ZN(\U4/Z_26 ) );
  NOR2_X2 U340 ( .A1(\top_add/A[12] ), .A2(n584), .ZN(n585) );
  XNOR2_X2 U341 ( .A(n585), .B(\top_add/A[13] ), .ZN(n586) );
  NOR2_X2 U342 ( .A1(n587), .A2(n586), .ZN(\U4/Z_27 ) );
  XOR2_X2 U343 ( .A(\bottom_add/A[8] ), .B(n18), .Z(n588) );
  NOR2_X2 U344 ( .A1(n588), .A2(n600), .ZN(\U6/Z_1 ) );
  NAND2_X2 U345 ( .A1(n18), .A2(n311), .ZN(n589) );
  XOR2_X2 U346 ( .A(n589), .B(n17), .Z(n590) );
  NOR2_X2 U347 ( .A1(n600), .A2(n590), .ZN(\U6/Z_2 ) );
  XOR2_X2 U348 ( .A(n591), .B(n16), .Z(n592) );
  NOR2_X2 U349 ( .A1(n600), .A2(n592), .ZN(\U6/Z_3 ) );
  NAND2_X2 U350 ( .A1(n593), .A2(n16), .ZN(n594) );
  XOR2_X2 U351 ( .A(n594), .B(n15), .Z(n595) );
  NOR2_X2 U352 ( .A1(n600), .A2(n595), .ZN(\U6/Z_4 ) );
  XOR2_X2 U353 ( .A(n596), .B(n14), .Z(n597) );
  NOR2_X2 U354 ( .A1(n600), .A2(n597), .ZN(\U6/Z_5 ) );
  NAND2_X2 U355 ( .A1(n14), .A2(n598), .ZN(n599) );
  XOR2_X2 U356 ( .A(n599), .B(n13), .Z(n601) );
  NOR2_X2 U357 ( .A1(n601), .A2(n600), .ZN(\U6/Z_6 ) );
  AND2_X1 U358 ( .A1(\U4/DATA1_0 ), .A2(n81), .ZN(\U4/Z_0 ) );
endmodule


module divider_pipe_stage_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n47, n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n62, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n85, n87, n88, n89, n90, n91, n92, n95, n96, n97,
         n98, n100, n102, n103, n104, n105, n106, n107, n108, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n128, n130, n131, n133, n134, n135, n139, n141,
         n145, n146, n147, n148, n149, n218, n219, n220, n221, n222, n223;

  XNOR2_X2 U2 ( .A(n29), .B(n3), .ZN(SUM[19]) );
  NAND2_X2 U4 ( .A1(n32), .A2(n25), .ZN(n23) );
  AOI21_X4 U5 ( .B1(n33), .B2(n25), .A(n26), .ZN(n24) );
  XNOR2_X2 U12 ( .A(n36), .B(n4), .ZN(SUM[18]) );
  NAND2_X2 U18 ( .A1(n133), .A2(n35), .ZN(n4) );
  NAND2_X2 U21 ( .A1(B[18]), .A2(A[18]), .ZN(n35) );
  NAND2_X2 U24 ( .A1(n134), .A2(n38), .ZN(n5) );
  NAND2_X2 U27 ( .A1(B[17]), .A2(A[17]), .ZN(n38) );
  XNOR2_X2 U28 ( .A(n43), .B(n6), .ZN(SUM[16]) );
  NAND2_X2 U32 ( .A1(n135), .A2(n42), .ZN(n6) );
  NAND2_X2 U35 ( .A1(B[16]), .A2(A[16]), .ZN(n42) );
  XNOR2_X2 U36 ( .A(n50), .B(n7), .ZN(SUM[15]) );
  NAND2_X2 U38 ( .A1(n219), .A2(n53), .ZN(n44) );
  NAND2_X2 U45 ( .A1(B[15]), .A2(A[15]), .ZN(n49) );
  XOR2_X2 U46 ( .A(n8), .B(n57), .Z(SUM[14]) );
  NAND2_X2 U52 ( .A1(n53), .A2(n52), .ZN(n8) );
  NAND2_X2 U55 ( .A1(B[14]), .A2(A[14]), .ZN(n52) );
  XOR2_X2 U56 ( .A(n9), .B(n65), .Z(SUM[13]) );
  NAND2_X2 U59 ( .A1(n66), .A2(n222), .ZN(n59) );
  NAND2_X2 U63 ( .A1(n222), .A2(n64), .ZN(n9) );
  NAND2_X2 U66 ( .A1(B[13]), .A2(A[13]), .ZN(n64) );
  XOR2_X2 U67 ( .A(n10), .B(n70), .Z(SUM[12]) );
  NAND2_X2 U71 ( .A1(n139), .A2(n69), .ZN(n10) );
  NAND2_X2 U74 ( .A1(B[12]), .A2(A[12]), .ZN(n69) );
  XNOR2_X2 U75 ( .A(n75), .B(n11), .ZN(SUM[11]) );
  NAND2_X2 U79 ( .A1(n71), .A2(n74), .ZN(n11) );
  NAND2_X2 U82 ( .A1(B[11]), .A2(A[11]), .ZN(n74) );
  XNOR2_X2 U83 ( .A(n81), .B(n12), .ZN(SUM[10]) );
  NAND2_X2 U88 ( .A1(n141), .A2(n80), .ZN(n12) );
  NAND2_X2 U91 ( .A1(B[10]), .A2(A[10]), .ZN(n80) );
  XNOR2_X2 U92 ( .A(n88), .B(n13), .ZN(SUM[9]) );
  NAND2_X2 U94 ( .A1(n220), .A2(n91), .ZN(n82) );
  NAND2_X2 U98 ( .A1(n220), .A2(n87), .ZN(n13) );
  NAND2_X2 U101 ( .A1(B[9]), .A2(A[9]), .ZN(n87) );
  XOR2_X2 U102 ( .A(n14), .B(n95), .Z(SUM[8]) );
  NAND2_X2 U108 ( .A1(n91), .A2(n90), .ZN(n14) );
  NAND2_X2 U111 ( .A1(B[8]), .A2(A[8]), .ZN(n90) );
  XOR2_X2 U112 ( .A(n15), .B(n103), .Z(SUM[7]) );
  NAND2_X2 U115 ( .A1(n104), .A2(n221), .ZN(n97) );
  NAND2_X2 U119 ( .A1(n221), .A2(n102), .ZN(n15) );
  NAND2_X2 U122 ( .A1(B[7]), .A2(A[7]), .ZN(n102) );
  XOR2_X2 U123 ( .A(n16), .B(n108), .Z(SUM[6]) );
  NAND2_X2 U127 ( .A1(n145), .A2(n107), .ZN(n16) );
  NAND2_X2 U130 ( .A1(B[6]), .A2(A[6]), .ZN(n107) );
  XNOR2_X2 U131 ( .A(n113), .B(n17), .ZN(SUM[5]) );
  NAND2_X2 U135 ( .A1(n146), .A2(n112), .ZN(n17) );
  NAND2_X2 U138 ( .A1(B[5]), .A2(A[5]), .ZN(n112) );
  XNOR2_X2 U139 ( .A(n119), .B(n18), .ZN(SUM[4]) );
  NAND2_X2 U144 ( .A1(n147), .A2(n118), .ZN(n18) );
  NAND2_X2 U147 ( .A1(B[4]), .A2(A[4]), .ZN(n118) );
  XOR2_X2 U148 ( .A(n19), .B(n122), .Z(SUM[3]) );
  NAND2_X2 U150 ( .A1(n148), .A2(n121), .ZN(n19) );
  NAND2_X2 U153 ( .A1(B[3]), .A2(A[3]), .ZN(n121) );
  XOR2_X2 U154 ( .A(n20), .B(n126), .Z(SUM[2]) );
  NAND2_X2 U157 ( .A1(n149), .A2(n125), .ZN(n20) );
  NAND2_X2 U160 ( .A1(B[2]), .A2(A[2]), .ZN(n125) );
  XOR2_X2 U161 ( .A(n131), .B(n21), .Z(SUM[1]) );
  NAND2_X2 U166 ( .A1(n223), .A2(n130), .ZN(n21) );
  NAND2_X2 U169 ( .A1(B[1]), .A2(A[1]), .ZN(n130) );
  XNOR2_X2 U170 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  AOI21_X2 U175 ( .B1(n58), .B2(n39), .A(n40), .ZN(n218) );
  AOI21_X2 U176 ( .B1(n58), .B2(n39), .A(n40), .ZN(n1) );
  NOR2_X2 U177 ( .A1(B[16]), .A2(A[16]), .ZN(n41) );
  AOI21_X2 U178 ( .B1(n219), .B2(n54), .A(n47), .ZN(n45) );
  NAND2_X2 U179 ( .A1(B[19]), .A2(A[19]), .ZN(n28) );
  AOI21_X2 U180 ( .B1(n96), .B2(n77), .A(n78), .ZN(n76) );
  OAI21_X2 U181 ( .B1(n76), .B2(n59), .A(n60), .ZN(n58) );
  INV_X2 U182 ( .A(n49), .ZN(n47) );
  NAND2_X1 U183 ( .A1(n219), .A2(n49), .ZN(n7) );
  INV_X4 U184 ( .A(n28), .ZN(n26) );
  XOR2_X1 U185 ( .A(n5), .B(n218), .Z(SUM[17]) );
  NAND2_X1 U186 ( .A1(n25), .A2(n28), .ZN(n3) );
  OAI21_X2 U187 ( .B1(n34), .B2(n38), .A(n35), .ZN(n33) );
  OR2_X2 U188 ( .A1(B[15]), .A2(A[15]), .ZN(n219) );
  OAI21_X1 U189 ( .B1(n218), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X1 U190 ( .B1(n218), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X2 U191 ( .B1(n1), .B2(n23), .A(n24), .ZN(CO) );
  INV_X1 U192 ( .A(n33), .ZN(n31) );
  OAI21_X1 U193 ( .B1(n95), .B2(n82), .A(n83), .ZN(n81) );
  OAI21_X1 U194 ( .B1(n57), .B2(n44), .A(n45), .ZN(n43) );
  NOR2_X2 U195 ( .A1(n41), .A2(n44), .ZN(n39) );
  INV_X2 U196 ( .A(n87), .ZN(n85) );
  AOI21_X2 U197 ( .B1(n113), .B2(n104), .A(n105), .ZN(n103) );
  AOI21_X2 U198 ( .B1(n75), .B2(n66), .A(n67), .ZN(n65) );
  OAI21_X2 U199 ( .B1(n45), .B2(n41), .A(n42), .ZN(n40) );
  AOI21_X2 U200 ( .B1(n220), .B2(n92), .A(n85), .ZN(n83) );
  AOI21_X2 U201 ( .B1(n223), .B2(n2), .A(n128), .ZN(n126) );
  AOI21_X2 U202 ( .B1(n123), .B2(n115), .A(n116), .ZN(n114) );
  NOR2_X2 U203 ( .A1(n117), .A2(n120), .ZN(n115) );
  OAI21_X2 U204 ( .B1(n117), .B2(n121), .A(n118), .ZN(n116) );
  NOR2_X2 U205 ( .A1(n82), .A2(n79), .ZN(n77) );
  OAI21_X2 U206 ( .B1(n83), .B2(n79), .A(n80), .ZN(n78) );
  OAI21_X2 U207 ( .B1(n106), .B2(n112), .A(n107), .ZN(n105) );
  OAI21_X2 U208 ( .B1(n68), .B2(n74), .A(n69), .ZN(n67) );
  OAI21_X2 U209 ( .B1(n126), .B2(n124), .A(n125), .ZN(n123) );
  AOI21_X2 U210 ( .B1(n67), .B2(n222), .A(n62), .ZN(n60) );
  OAI21_X2 U211 ( .B1(n114), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X2 U212 ( .B1(n105), .B2(n221), .A(n100), .ZN(n98) );
  AOI21_X2 U213 ( .B1(n113), .B2(n146), .A(n110), .ZN(n108) );
  AOI21_X2 U214 ( .B1(n75), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U215 ( .B1(n95), .B2(n89), .A(n90), .ZN(n88) );
  OAI21_X1 U216 ( .B1(n57), .B2(n51), .A(n52), .ZN(n50) );
  NOR2_X2 U217 ( .A1(n106), .A2(n111), .ZN(n104) );
  NOR2_X2 U218 ( .A1(n68), .A2(n73), .ZN(n66) );
  NOR2_X2 U219 ( .A1(n34), .A2(n37), .ZN(n32) );
  OAI21_X2 U220 ( .B1(n122), .B2(n120), .A(n121), .ZN(n119) );
  NOR2_X2 U221 ( .A1(B[17]), .A2(A[17]), .ZN(n37) );
  NOR2_X2 U222 ( .A1(B[10]), .A2(A[10]), .ZN(n79) );
  NOR2_X2 U223 ( .A1(B[3]), .A2(A[3]), .ZN(n120) );
  NOR2_X2 U224 ( .A1(B[18]), .A2(A[18]), .ZN(n34) );
  NOR2_X2 U225 ( .A1(B[6]), .A2(A[6]), .ZN(n106) );
  NOR2_X2 U226 ( .A1(B[12]), .A2(A[12]), .ZN(n68) );
  NOR2_X2 U227 ( .A1(B[4]), .A2(A[4]), .ZN(n117) );
  NOR2_X2 U228 ( .A1(B[5]), .A2(A[5]), .ZN(n111) );
  NOR2_X2 U229 ( .A1(B[11]), .A2(A[11]), .ZN(n73) );
  NOR2_X1 U230 ( .A1(B[8]), .A2(A[8]), .ZN(n89) );
  NOR2_X1 U231 ( .A1(B[14]), .A2(A[14]), .ZN(n51) );
  NOR2_X2 U232 ( .A1(B[2]), .A2(A[2]), .ZN(n124) );
  NOR2_X2 U233 ( .A1(B[0]), .A2(A[0]), .ZN(n131) );
  OR2_X1 U234 ( .A1(B[9]), .A2(A[9]), .ZN(n220) );
  NOR2_X2 U235 ( .A1(B[19]), .A2(A[19]), .ZN(n27) );
  OR2_X1 U236 ( .A1(B[7]), .A2(A[7]), .ZN(n221) );
  OR2_X1 U237 ( .A1(B[13]), .A2(A[13]), .ZN(n222) );
  OR2_X1 U238 ( .A1(B[1]), .A2(A[1]), .ZN(n223) );
  INV_X4 U239 ( .A(n96), .ZN(n95) );
  INV_X4 U240 ( .A(n90), .ZN(n92) );
  INV_X4 U241 ( .A(n76), .ZN(n75) );
  INV_X4 U242 ( .A(n74), .ZN(n72) );
  INV_X4 U243 ( .A(n64), .ZN(n62) );
  INV_X4 U244 ( .A(n58), .ZN(n57) );
  INV_X4 U245 ( .A(n52), .ZN(n54) );
  INV_X4 U246 ( .A(n32), .ZN(n30) );
  INV_X4 U247 ( .A(n131), .ZN(n2) );
  INV_X4 U248 ( .A(n124), .ZN(n149) );
  INV_X4 U249 ( .A(n120), .ZN(n148) );
  INV_X4 U250 ( .A(n117), .ZN(n147) );
  INV_X4 U251 ( .A(n106), .ZN(n145) );
  INV_X4 U252 ( .A(n89), .ZN(n91) );
  INV_X4 U253 ( .A(n79), .ZN(n141) );
  INV_X4 U254 ( .A(n73), .ZN(n71) );
  INV_X4 U255 ( .A(n68), .ZN(n139) );
  INV_X4 U256 ( .A(n51), .ZN(n53) );
  INV_X4 U257 ( .A(n41), .ZN(n135) );
  INV_X4 U258 ( .A(n37), .ZN(n134) );
  INV_X4 U259 ( .A(n34), .ZN(n133) );
  INV_X4 U260 ( .A(n27), .ZN(n25) );
  INV_X4 U261 ( .A(n130), .ZN(n128) );
  INV_X4 U262 ( .A(n123), .ZN(n122) );
  INV_X4 U263 ( .A(n114), .ZN(n113) );
  INV_X4 U264 ( .A(n112), .ZN(n110) );
  INV_X4 U265 ( .A(n111), .ZN(n146) );
  INV_X4 U266 ( .A(n102), .ZN(n100) );
endmodule


module divider_pipe_stage_1 ( clock, reset_n, start, divided, divisor, q_in, 
        start_out, divisor_out, result, q_out );
  input [27:0] divided;
  input [19:0] divisor;
  input [7:0] q_in;
  output [19:0] divisor_out;
  output [27:0] result;
  output [7:0] q_out;
  input clock, reset_n, start;
  output start_out;
  wire   N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N75,
         N76, N77, N78, N79, N80, N81, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319;
  wire   [20:0] stage_result;

  DFFR_X1 \q_out_reg[7]  ( .D(N81), .CK(clock), .RN(n233), .Q(q_out[7]) );
  DFFR_X1 \q_out_reg[6]  ( .D(N80), .CK(clock), .RN(n233), .Q(q_out[6]) );
  DFFR_X1 \q_out_reg[5]  ( .D(N79), .CK(clock), .RN(n233), .Q(q_out[5]) );
  DFFR_X1 \q_out_reg[4]  ( .D(N78), .CK(clock), .RN(n233), .Q(q_out[4]) );
  DFFR_X1 \q_out_reg[3]  ( .D(N77), .CK(clock), .RN(n233), .Q(q_out[3]) );
  DFFR_X1 \q_out_reg[2]  ( .D(N76), .CK(clock), .RN(n233), .Q(q_out[2]) );
  DFFR_X1 \q_out_reg[1]  ( .D(N75), .CK(clock), .RN(n233), .Q(q_out[1]) );
  DFFR_X1 \divisor_out_reg[19]  ( .D(N46), .CK(clock), .RN(n230), .Q(
        divisor_out[19]) );
  DFFR_X1 \divisor_out_reg[18]  ( .D(N45), .CK(clock), .RN(n233), .Q(
        divisor_out[18]) );
  DFFR_X1 \divisor_out_reg[17]  ( .D(N44), .CK(clock), .RN(n232), .Q(
        divisor_out[17]) );
  DFFR_X1 \divisor_out_reg[16]  ( .D(N43), .CK(clock), .RN(n231), .Q(
        divisor_out[16]) );
  DFFR_X1 \divisor_out_reg[15]  ( .D(N42), .CK(clock), .RN(n233), .Q(
        divisor_out[15]) );
  DFFR_X1 \divisor_out_reg[14]  ( .D(N41), .CK(clock), .RN(n232), .Q(
        divisor_out[14]) );
  DFFR_X1 \divisor_out_reg[13]  ( .D(N40), .CK(clock), .RN(n231), .Q(
        divisor_out[13]) );
  DFFR_X1 \divisor_out_reg[12]  ( .D(N39), .CK(clock), .RN(n233), .Q(
        divisor_out[12]) );
  DFFR_X1 \divisor_out_reg[11]  ( .D(N38), .CK(clock), .RN(n230), .Q(
        divisor_out[11]) );
  DFFR_X1 \divisor_out_reg[10]  ( .D(N37), .CK(clock), .RN(n230), .Q(
        divisor_out[10]) );
  DFFR_X1 \divisor_out_reg[9]  ( .D(N36), .CK(clock), .RN(n230), .Q(
        divisor_out[9]) );
  DFFR_X1 \divisor_out_reg[8]  ( .D(N35), .CK(clock), .RN(n230), .Q(
        divisor_out[8]) );
  DFFR_X1 \divisor_out_reg[7]  ( .D(N34), .CK(clock), .RN(n230), .Q(
        divisor_out[7]) );
  DFFR_X1 \divisor_out_reg[6]  ( .D(N33), .CK(clock), .RN(n230), .Q(
        divisor_out[6]) );
  DFFR_X1 \divisor_out_reg[5]  ( .D(N32), .CK(clock), .RN(n230), .Q(
        divisor_out[5]) );
  DFFR_X1 \divisor_out_reg[4]  ( .D(N31), .CK(clock), .RN(n230), .Q(
        divisor_out[4]) );
  DFFR_X1 \divisor_out_reg[3]  ( .D(N30), .CK(clock), .RN(n230), .Q(
        divisor_out[3]) );
  DFFR_X1 \divisor_out_reg[2]  ( .D(N29), .CK(clock), .RN(n230), .Q(
        divisor_out[2]) );
  DFFR_X1 \divisor_out_reg[1]  ( .D(N28), .CK(clock), .RN(n230), .Q(
        divisor_out[1]) );
  DFFR_X1 \divisor_out_reg[0]  ( .D(N27), .CK(clock), .RN(n230), .Q(
        divisor_out[0]) );
  AND2_X1 U47 ( .A1(start), .A2(q_in[6]), .ZN(N81) );
  AND2_X1 U48 ( .A1(q_in[5]), .A2(start), .ZN(N80) );
  AND2_X1 U49 ( .A1(q_in[4]), .A2(start), .ZN(N79) );
  AND2_X1 U50 ( .A1(q_in[3]), .A2(start), .ZN(N78) );
  AND2_X1 U51 ( .A1(q_in[2]), .A2(start), .ZN(N77) );
  AND2_X1 U52 ( .A1(q_in[1]), .A2(start), .ZN(N76) );
  AND2_X1 U53 ( .A1(q_in[0]), .A2(start), .ZN(N75) );
  AND2_X1 U56 ( .A1(divided[5]), .A2(start), .ZN(N52) );
  AND2_X1 U57 ( .A1(divided[4]), .A2(start), .ZN(N51) );
  AND2_X1 U58 ( .A1(divided[3]), .A2(start), .ZN(N50) );
  AND2_X1 U59 ( .A1(divided[2]), .A2(start), .ZN(N49) );
  AND2_X1 U60 ( .A1(divided[1]), .A2(start), .ZN(N48) );
  AND2_X1 U61 ( .A1(divided[0]), .A2(start), .ZN(N47) );
  divider_pipe_stage_1_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  DFFR_X1 \result_reg[27]  ( .D(n319), .CK(clock), .RN(n232), .Q(result[27])
         );
  DFFR_X1 \result_reg[23]  ( .D(n315), .CK(clock), .RN(n232), .Q(result[23])
         );
  DFFR_X1 \result_reg[25]  ( .D(n317), .CK(clock), .RN(n232), .Q(result[25])
         );
  DFFR_X1 \result_reg[8]  ( .D(n300), .CK(clock), .RN(n231), .Q(result[8]) );
  DFFR_X1 \result_reg[13]  ( .D(n305), .CK(clock), .RN(n231), .Q(result[13])
         );
  DFFR_X1 \result_reg[11]  ( .D(n303), .CK(clock), .RN(n231), .Q(result[11])
         );
  DFFR_X1 \result_reg[9]  ( .D(n301), .CK(clock), .RN(n231), .Q(result[9]) );
  DFFR_X1 \result_reg[19]  ( .D(n311), .CK(clock), .RN(n232), .Q(result[19])
         );
  DFFR_X1 \result_reg[15]  ( .D(n307), .CK(clock), .RN(n231), .Q(result[15])
         );
  DFFR_X1 \result_reg[21]  ( .D(n313), .CK(clock), .RN(n232), .Q(result[21])
         );
  DFFR_X1 \result_reg[17]  ( .D(n309), .CK(clock), .RN(n232), .Q(result[17])
         );
  DFFR_X2 start_out_reg ( .D(start), .CK(clock), .RN(n233), .Q(start_out) );
  DFFR_X2 \result_reg[7]  ( .D(N53), .CK(clock), .RN(n231), .Q(result[7]) );
  DFFR_X2 \result_reg[6]  ( .D(N52), .CK(clock), .RN(n231), .Q(result[6]) );
  DFFR_X2 \result_reg[5]  ( .D(N51), .CK(clock), .RN(n231), .Q(result[5]) );
  DFFR_X2 \result_reg[4]  ( .D(N50), .CK(clock), .RN(n233), .Q(result[4]) );
  DFFR_X2 \result_reg[3]  ( .D(N49), .CK(clock), .RN(n230), .Q(result[3]) );
  DFFR_X2 \result_reg[2]  ( .D(N48), .CK(clock), .RN(n233), .Q(result[2]) );
  DFFR_X2 \result_reg[1]  ( .D(N47), .CK(clock), .RN(n233), .Q(result[1]) );
  DFFR_X2 \q_out_reg[0]  ( .D(n299), .CK(clock), .RN(n232), .Q(q_out[0]) );
  DFFR_X2 \result_reg[24]  ( .D(n316), .CK(clock), .RN(n232), .Q(result[24])
         );
  DFFR_X2 \result_reg[26]  ( .D(n318), .CK(clock), .RN(n232), .Q(result[26])
         );
  DFFR_X2 \result_reg[20]  ( .D(n312), .CK(clock), .RN(n232), .Q(result[20])
         );
  DFFR_X2 \result_reg[18]  ( .D(n310), .CK(clock), .RN(n232), .Q(result[18])
         );
  DFFR_X2 \result_reg[14]  ( .D(n306), .CK(clock), .RN(n231), .Q(result[14])
         );
  DFFR_X2 \result_reg[12]  ( .D(n304), .CK(clock), .RN(n231), .Q(result[12])
         );
  DFFR_X2 \result_reg[10]  ( .D(n302), .CK(clock), .RN(n231), .Q(result[10])
         );
  DFFR_X2 \result_reg[22]  ( .D(n314), .CK(clock), .RN(n232), .Q(result[22])
         );
  DFFR_X2 \result_reg[16]  ( .D(n308), .CK(clock), .RN(n231), .Q(result[16])
         );
  INV_X4 U4 ( .A(1'b1), .ZN(result[0]) );
  INV_X16 U6 ( .A(n227), .ZN(n229) );
  INV_X16 U7 ( .A(n225), .ZN(n226) );
  AND2_X4 U8 ( .A1(start), .A2(n236), .ZN(n225) );
  AND2_X4 U9 ( .A1(start), .A2(n236), .ZN(n227) );
  INV_X1 U10 ( .A(divisor[19]), .ZN(n297) );
  INV_X4 U11 ( .A(n234), .ZN(n231) );
  INV_X4 U12 ( .A(n234), .ZN(n232) );
  INV_X4 U13 ( .A(n234), .ZN(n230) );
  INV_X4 U14 ( .A(n234), .ZN(n233) );
  INV_X4 U15 ( .A(reset_n), .ZN(n234) );
  INV_X2 U16 ( .A(start), .ZN(n298) );
  NAND2_X4 U17 ( .A1(start), .A2(n235), .ZN(n228) );
  NAND2_X4 U18 ( .A1(start), .A2(n235), .ZN(n276) );
  XNOR2_X2 U19 ( .A(divided[27]), .B(stage_result[20]), .ZN(n236) );
  INV_X4 U20 ( .A(n236), .ZN(n235) );
  INV_X4 U21 ( .A(n276), .ZN(n299) );
  AND2_X1 U22 ( .A1(divided[6]), .A2(start), .ZN(N53) );
  INV_X4 U23 ( .A(divided[7]), .ZN(n238) );
  INV_X4 U24 ( .A(stage_result[0]), .ZN(n237) );
  OAI22_X2 U25 ( .A1(n229), .A2(n238), .B1(n228), .B2(n237), .ZN(n300) );
  INV_X4 U26 ( .A(divided[8]), .ZN(n240) );
  INV_X4 U27 ( .A(stage_result[1]), .ZN(n239) );
  OAI22_X2 U28 ( .A1(n226), .A2(n240), .B1(n228), .B2(n239), .ZN(n301) );
  INV_X4 U29 ( .A(divided[9]), .ZN(n242) );
  INV_X4 U30 ( .A(stage_result[2]), .ZN(n241) );
  OAI22_X2 U31 ( .A1(n229), .A2(n242), .B1(n276), .B2(n241), .ZN(n302) );
  INV_X4 U32 ( .A(divided[10]), .ZN(n244) );
  INV_X4 U33 ( .A(stage_result[3]), .ZN(n243) );
  OAI22_X2 U34 ( .A1(n226), .A2(n244), .B1(n228), .B2(n243), .ZN(n303) );
  INV_X4 U35 ( .A(divided[11]), .ZN(n246) );
  INV_X4 U36 ( .A(stage_result[4]), .ZN(n245) );
  OAI22_X2 U37 ( .A1(n229), .A2(n246), .B1(n276), .B2(n245), .ZN(n304) );
  INV_X4 U38 ( .A(divided[12]), .ZN(n248) );
  INV_X4 U39 ( .A(stage_result[5]), .ZN(n247) );
  OAI22_X2 U40 ( .A1(n226), .A2(n248), .B1(n228), .B2(n247), .ZN(n305) );
  INV_X4 U41 ( .A(divided[13]), .ZN(n250) );
  INV_X4 U42 ( .A(stage_result[6]), .ZN(n249) );
  OAI22_X2 U43 ( .A1(n229), .A2(n250), .B1(n276), .B2(n249), .ZN(n306) );
  INV_X4 U44 ( .A(divided[14]), .ZN(n252) );
  INV_X4 U45 ( .A(stage_result[7]), .ZN(n251) );
  OAI22_X2 U46 ( .A1(n226), .A2(n252), .B1(n228), .B2(n251), .ZN(n307) );
  INV_X4 U54 ( .A(divided[15]), .ZN(n254) );
  INV_X4 U55 ( .A(stage_result[8]), .ZN(n253) );
  OAI22_X2 U62 ( .A1(n229), .A2(n254), .B1(n276), .B2(n253), .ZN(n308) );
  INV_X4 U63 ( .A(divided[16]), .ZN(n256) );
  INV_X4 U64 ( .A(stage_result[9]), .ZN(n255) );
  OAI22_X2 U65 ( .A1(n226), .A2(n256), .B1(n228), .B2(n255), .ZN(n309) );
  INV_X4 U66 ( .A(divided[17]), .ZN(n258) );
  INV_X4 U67 ( .A(stage_result[10]), .ZN(n257) );
  OAI22_X2 U68 ( .A1(n229), .A2(n258), .B1(n276), .B2(n257), .ZN(n310) );
  INV_X4 U69 ( .A(divided[18]), .ZN(n260) );
  INV_X4 U70 ( .A(stage_result[11]), .ZN(n259) );
  OAI22_X2 U71 ( .A1(n226), .A2(n260), .B1(n228), .B2(n259), .ZN(n311) );
  INV_X4 U72 ( .A(divided[19]), .ZN(n262) );
  INV_X4 U73 ( .A(stage_result[12]), .ZN(n261) );
  OAI22_X2 U74 ( .A1(n229), .A2(n262), .B1(n276), .B2(n261), .ZN(n312) );
  INV_X4 U75 ( .A(divided[20]), .ZN(n264) );
  INV_X4 U76 ( .A(stage_result[13]), .ZN(n263) );
  OAI22_X2 U77 ( .A1(n226), .A2(n264), .B1(n228), .B2(n263), .ZN(n313) );
  INV_X4 U78 ( .A(divided[21]), .ZN(n266) );
  INV_X4 U79 ( .A(stage_result[14]), .ZN(n265) );
  OAI22_X2 U80 ( .A1(n229), .A2(n266), .B1(n276), .B2(n265), .ZN(n314) );
  INV_X4 U81 ( .A(divided[22]), .ZN(n268) );
  INV_X4 U82 ( .A(stage_result[15]), .ZN(n267) );
  OAI22_X2 U83 ( .A1(n226), .A2(n268), .B1(n228), .B2(n267), .ZN(n315) );
  INV_X4 U84 ( .A(divided[23]), .ZN(n270) );
  INV_X4 U85 ( .A(stage_result[16]), .ZN(n269) );
  OAI22_X2 U86 ( .A1(n229), .A2(n270), .B1(n276), .B2(n269), .ZN(n316) );
  INV_X4 U87 ( .A(divided[24]), .ZN(n272) );
  INV_X4 U88 ( .A(stage_result[17]), .ZN(n271) );
  OAI22_X2 U89 ( .A1(n226), .A2(n272), .B1(n228), .B2(n271), .ZN(n317) );
  INV_X4 U90 ( .A(divided[25]), .ZN(n274) );
  INV_X4 U91 ( .A(stage_result[18]), .ZN(n273) );
  OAI22_X2 U92 ( .A1(n229), .A2(n274), .B1(n276), .B2(n273), .ZN(n318) );
  INV_X4 U93 ( .A(divided[26]), .ZN(n277) );
  INV_X4 U94 ( .A(stage_result[19]), .ZN(n275) );
  OAI22_X2 U95 ( .A1(n226), .A2(n277), .B1(n228), .B2(n275), .ZN(n319) );
  INV_X4 U96 ( .A(divisor[0]), .ZN(n278) );
  NOR2_X2 U97 ( .A1(n298), .A2(n278), .ZN(N27) );
  INV_X4 U98 ( .A(divisor[1]), .ZN(n279) );
  NOR2_X2 U99 ( .A1(n298), .A2(n279), .ZN(N28) );
  INV_X4 U100 ( .A(divisor[2]), .ZN(n280) );
  NOR2_X2 U101 ( .A1(n298), .A2(n280), .ZN(N29) );
  INV_X4 U102 ( .A(divisor[3]), .ZN(n281) );
  NOR2_X2 U103 ( .A1(n298), .A2(n281), .ZN(N30) );
  INV_X4 U104 ( .A(divisor[4]), .ZN(n282) );
  NOR2_X2 U105 ( .A1(n298), .A2(n282), .ZN(N31) );
  INV_X4 U106 ( .A(divisor[5]), .ZN(n283) );
  NOR2_X2 U107 ( .A1(n298), .A2(n283), .ZN(N32) );
  INV_X4 U108 ( .A(divisor[6]), .ZN(n284) );
  NOR2_X2 U109 ( .A1(n298), .A2(n284), .ZN(N33) );
  INV_X4 U110 ( .A(divisor[7]), .ZN(n285) );
  NOR2_X2 U111 ( .A1(n298), .A2(n285), .ZN(N34) );
  INV_X4 U112 ( .A(divisor[8]), .ZN(n286) );
  NOR2_X2 U113 ( .A1(n298), .A2(n286), .ZN(N35) );
  INV_X4 U114 ( .A(divisor[9]), .ZN(n287) );
  NOR2_X2 U115 ( .A1(n298), .A2(n287), .ZN(N36) );
  INV_X4 U116 ( .A(divisor[10]), .ZN(n288) );
  NOR2_X2 U117 ( .A1(n298), .A2(n288), .ZN(N37) );
  INV_X4 U118 ( .A(divisor[11]), .ZN(n289) );
  NOR2_X2 U119 ( .A1(n298), .A2(n289), .ZN(N38) );
  INV_X4 U120 ( .A(divisor[12]), .ZN(n290) );
  NOR2_X2 U121 ( .A1(n298), .A2(n290), .ZN(N39) );
  INV_X4 U122 ( .A(divisor[13]), .ZN(n291) );
  NOR2_X2 U123 ( .A1(n298), .A2(n291), .ZN(N40) );
  INV_X4 U124 ( .A(divisor[14]), .ZN(n292) );
  NOR2_X2 U125 ( .A1(n298), .A2(n292), .ZN(N41) );
  INV_X4 U126 ( .A(divisor[15]), .ZN(n293) );
  NOR2_X2 U127 ( .A1(n298), .A2(n293), .ZN(N42) );
  INV_X4 U128 ( .A(divisor[16]), .ZN(n294) );
  NOR2_X2 U129 ( .A1(n298), .A2(n294), .ZN(N43) );
  INV_X4 U130 ( .A(divisor[17]), .ZN(n295) );
  NOR2_X2 U131 ( .A1(n298), .A2(n295), .ZN(N44) );
  INV_X4 U132 ( .A(divisor[18]), .ZN(n296) );
  NOR2_X2 U133 ( .A1(n298), .A2(n296), .ZN(N45) );
  NOR2_X2 U134 ( .A1(n298), .A2(n297), .ZN(N46) );
endmodule


module divider_pipe_stage_6_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n110, n112, n114,
         n115, n116, n117, n118, n120, n121, n122;

  FA_X1 U2 ( .A(A[19]), .B(B[19]), .CI(n18), .CO(CO), .S(SUM[19]) );
  FA_X1 U3 ( .A(A[18]), .B(B[18]), .CI(n19), .CO(n18), .S(SUM[18]) );
  FA_X1 U4 ( .A(A[17]), .B(B[17]), .CI(n20), .CO(n19), .S(SUM[17]) );
  XOR2_X2 U5 ( .A(n1), .B(n23), .Z(SUM[16]) );
  NAND2_X2 U7 ( .A1(n107), .A2(n22), .ZN(n1) );
  NAND2_X2 U10 ( .A1(A[16]), .A2(B[16]), .ZN(n22) );
  XOR2_X2 U11 ( .A(n2), .B(n32), .Z(SUM[15]) );
  NAND2_X2 U15 ( .A1(n40), .A2(n28), .ZN(n26) );
  NAND2_X2 U19 ( .A1(n108), .A2(n31), .ZN(n2) );
  NAND2_X2 U22 ( .A1(A[15]), .A2(B[15]), .ZN(n31) );
  XNOR2_X2 U23 ( .A(n37), .B(n3), .ZN(SUM[14]) );
  NAND2_X2 U27 ( .A1(n33), .A2(n36), .ZN(n3) );
  NAND2_X2 U30 ( .A1(A[14]), .A2(B[14]), .ZN(n36) );
  XOR2_X2 U31 ( .A(n4), .B(n44), .Z(SUM[13]) );
  NAND2_X2 U37 ( .A1(n110), .A2(n43), .ZN(n4) );
  NAND2_X2 U40 ( .A1(A[13]), .A2(B[13]), .ZN(n43) );
  XOR2_X2 U41 ( .A(n5), .B(n49), .Z(SUM[12]) );
  NAND2_X2 U45 ( .A1(n45), .A2(n48), .ZN(n5) );
  NAND2_X2 U48 ( .A1(A[12]), .A2(B[12]), .ZN(n48) );
  XOR2_X2 U49 ( .A(n6), .B(n57), .Z(SUM[11]) );
  NAND2_X2 U52 ( .A1(n65), .A2(n53), .ZN(n51) );
  NAND2_X2 U56 ( .A1(n112), .A2(n56), .ZN(n6) );
  NAND2_X2 U59 ( .A1(A[11]), .A2(B[11]), .ZN(n56) );
  XNOR2_X2 U60 ( .A(n62), .B(n7), .ZN(SUM[10]) );
  NAND2_X2 U64 ( .A1(n58), .A2(n61), .ZN(n7) );
  NAND2_X2 U67 ( .A1(A[10]), .A2(B[10]), .ZN(n61) );
  XNOR2_X2 U68 ( .A(n69), .B(n8), .ZN(SUM[9]) );
  NAND2_X2 U74 ( .A1(n114), .A2(n68), .ZN(n8) );
  NAND2_X2 U77 ( .A1(A[9]), .A2(B[9]), .ZN(n68) );
  XOR2_X2 U78 ( .A(n9), .B(n72), .Z(SUM[8]) );
  NAND2_X2 U80 ( .A1(n115), .A2(n71), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[8]), .A2(B[8]), .ZN(n71) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[7]) );
  NAND2_X2 U87 ( .A1(n84), .A2(n76), .ZN(n74) );
  NAND2_X2 U91 ( .A1(n116), .A2(n79), .ZN(n10) );
  NAND2_X2 U94 ( .A1(A[7]), .A2(B[7]), .ZN(n79) );
  XOR2_X2 U95 ( .A(n11), .B(n83), .Z(SUM[6]) );
  NAND2_X2 U97 ( .A1(n117), .A2(n82), .ZN(n11) );
  NAND2_X2 U100 ( .A1(A[6]), .A2(B[6]), .ZN(n82) );
  XOR2_X2 U101 ( .A(n12), .B(n88), .Z(SUM[5]) );
  NAND2_X2 U105 ( .A1(n118), .A2(n87), .ZN(n12) );
  NAND2_X2 U108 ( .A1(A[5]), .A2(B[5]), .ZN(n87) );
  XNOR2_X2 U109 ( .A(n93), .B(n13), .ZN(SUM[4]) );
  NAND2_X2 U113 ( .A1(n89), .A2(n92), .ZN(n13) );
  NAND2_X2 U116 ( .A1(A[4]), .A2(B[4]), .ZN(n92) );
  XNOR2_X2 U117 ( .A(n99), .B(n14), .ZN(SUM[3]) );
  NAND2_X2 U122 ( .A1(n120), .A2(n98), .ZN(n14) );
  NAND2_X2 U125 ( .A1(A[3]), .A2(B[3]), .ZN(n98) );
  XOR2_X2 U126 ( .A(n15), .B(n102), .Z(SUM[2]) );
  NAND2_X2 U128 ( .A1(n121), .A2(n101), .ZN(n15) );
  NAND2_X2 U131 ( .A1(A[2]), .A2(B[2]), .ZN(n101) );
  XOR2_X2 U132 ( .A(n106), .B(n16), .Z(SUM[1]) );
  NAND2_X2 U135 ( .A1(n122), .A2(n105), .ZN(n16) );
  NAND2_X2 U138 ( .A1(A[1]), .A2(B[1]), .ZN(n105) );
  XNOR2_X2 U139 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U144 ( .B1(n73), .B2(n24), .A(n25), .ZN(n23) );
  NOR2_X2 U145 ( .A1(n51), .A2(n26), .ZN(n24) );
  OAI21_X2 U146 ( .B1(n52), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X2 U147 ( .B1(n49), .B2(n38), .A(n39), .ZN(n37) );
  OAI21_X2 U148 ( .B1(n72), .B2(n51), .A(n52), .ZN(n50) );
  AOI21_X2 U149 ( .B1(n93), .B2(n84), .A(n85), .ZN(n83) );
  OAI21_X2 U150 ( .B1(n72), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X2 U151 ( .B1(n53), .B2(n66), .A(n54), .ZN(n52) );
  OAI21_X2 U152 ( .B1(n55), .B2(n61), .A(n56), .ZN(n54) );
  AOI21_X2 U153 ( .B1(n95), .B2(n103), .A(n96), .ZN(n94) );
  NOR2_X2 U154 ( .A1(n100), .A2(n97), .ZN(n95) );
  OAI21_X2 U155 ( .B1(n97), .B2(n101), .A(n98), .ZN(n96) );
  OAI21_X2 U156 ( .B1(n86), .B2(n92), .A(n87), .ZN(n85) );
  OAI21_X2 U157 ( .B1(n94), .B2(n74), .A(n75), .ZN(n73) );
  AOI21_X2 U158 ( .B1(n76), .B2(n85), .A(n77), .ZN(n75) );
  NOR2_X2 U159 ( .A1(n81), .A2(n78), .ZN(n76) );
  AOI21_X2 U160 ( .B1(n28), .B2(n41), .A(n29), .ZN(n27) );
  OAI21_X2 U161 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  OAI21_X2 U162 ( .B1(n42), .B2(n48), .A(n43), .ZN(n41) );
  OAI21_X2 U163 ( .B1(n104), .B2(n106), .A(n105), .ZN(n103) );
  OAI21_X2 U164 ( .B1(n67), .B2(n71), .A(n68), .ZN(n66) );
  OAI21_X2 U165 ( .B1(n78), .B2(n82), .A(n79), .ZN(n77) );
  NOR2_X2 U166 ( .A1(n60), .A2(n55), .ZN(n53) );
  NOR2_X2 U167 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U168 ( .A1(n91), .A2(n86), .ZN(n84) );
  NOR2_X2 U169 ( .A1(n70), .A2(n67), .ZN(n65) );
  NOR2_X2 U170 ( .A1(n47), .A2(n42), .ZN(n40) );
  AOI21_X2 U171 ( .B1(n37), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U172 ( .B1(n93), .B2(n89), .A(n90), .ZN(n88) );
  AOI21_X2 U173 ( .B1(n62), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X2 U174 ( .B1(n50), .B2(n45), .A(n46), .ZN(n44) );
  OAI21_X2 U175 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X2 U176 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U177 ( .B1(n72), .B2(n70), .A(n71), .ZN(n69) );
  OAI21_X2 U178 ( .B1(n23), .B2(n21), .A(n22), .ZN(n20) );
  NOR2_X2 U179 ( .A1(A[3]), .A2(B[3]), .ZN(n97) );
  NOR2_X2 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n78) );
  NOR2_X2 U181 ( .A1(A[5]), .A2(B[5]), .ZN(n86) );
  NOR2_X2 U182 ( .A1(A[11]), .A2(B[11]), .ZN(n55) );
  NOR2_X2 U183 ( .A1(A[9]), .A2(B[9]), .ZN(n67) );
  NOR2_X2 U184 ( .A1(A[15]), .A2(B[15]), .ZN(n30) );
  NOR2_X2 U185 ( .A1(A[13]), .A2(B[13]), .ZN(n42) );
  NOR2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n100) );
  NOR2_X2 U187 ( .A1(A[6]), .A2(B[6]), .ZN(n81) );
  NOR2_X2 U188 ( .A1(A[8]), .A2(B[8]), .ZN(n70) );
  NOR2_X2 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n104) );
  NOR2_X2 U190 ( .A1(A[0]), .A2(B[0]), .ZN(n106) );
  NOR2_X2 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n91) );
  NOR2_X2 U192 ( .A1(A[10]), .A2(B[10]), .ZN(n60) );
  NOR2_X2 U193 ( .A1(A[12]), .A2(B[12]), .ZN(n47) );
  NOR2_X2 U194 ( .A1(A[14]), .A2(B[14]), .ZN(n35) );
  NOR2_X2 U195 ( .A1(A[16]), .A2(B[16]), .ZN(n21) );
  INV_X4 U196 ( .A(n94), .ZN(n93) );
  INV_X4 U197 ( .A(n92), .ZN(n90) );
  INV_X4 U198 ( .A(n73), .ZN(n72) );
  INV_X4 U199 ( .A(n66), .ZN(n64) );
  INV_X4 U200 ( .A(n65), .ZN(n63) );
  INV_X4 U201 ( .A(n61), .ZN(n59) );
  INV_X4 U202 ( .A(n50), .ZN(n49) );
  INV_X4 U203 ( .A(n48), .ZN(n46) );
  INV_X4 U204 ( .A(n41), .ZN(n39) );
  INV_X4 U205 ( .A(n40), .ZN(n38) );
  INV_X4 U206 ( .A(n36), .ZN(n34) );
  INV_X4 U207 ( .A(n104), .ZN(n122) );
  INV_X4 U208 ( .A(n100), .ZN(n121) );
  INV_X4 U209 ( .A(n97), .ZN(n120) );
  INV_X4 U210 ( .A(n91), .ZN(n89) );
  INV_X4 U211 ( .A(n86), .ZN(n118) );
  INV_X4 U212 ( .A(n81), .ZN(n117) );
  INV_X4 U213 ( .A(n78), .ZN(n116) );
  INV_X4 U214 ( .A(n70), .ZN(n115) );
  INV_X4 U215 ( .A(n67), .ZN(n114) );
  INV_X4 U216 ( .A(n60), .ZN(n58) );
  INV_X4 U217 ( .A(n55), .ZN(n112) );
  INV_X4 U218 ( .A(n47), .ZN(n45) );
  INV_X4 U219 ( .A(n42), .ZN(n110) );
  INV_X4 U220 ( .A(n35), .ZN(n33) );
  INV_X4 U221 ( .A(n30), .ZN(n108) );
  INV_X4 U222 ( .A(n21), .ZN(n107) );
  INV_X4 U223 ( .A(n103), .ZN(n102) );
endmodule


module divider_pipe_stage_6 ( clock, reset_n, start, divided, divisor, q_in, 
        start_out, divisor_out, result, q_out );
  input [27:0] divided;
  input [19:0] divisor;
  input [7:0] q_in;
  output [19:0] divisor_out;
  output [27:0] result;
  output [7:0] q_out;
  input clock, reset_n, start;
  output start_out;
  wire   N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N75,
         N76, N77, N78, N79, N80, N81, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312;
  wire   [20:0] stage_result;

  DFFR_X1 start_out_reg ( .D(start), .CK(clock), .RN(n233), .Q(start_out) );
  DFFR_X1 \q_out_reg[7]  ( .D(N81), .CK(clock), .RN(n233), .Q(q_out[7]) );
  DFFR_X1 \q_out_reg[6]  ( .D(N80), .CK(clock), .RN(n233), .Q(q_out[6]) );
  DFFR_X1 \q_out_reg[5]  ( .D(N79), .CK(clock), .RN(n233), .Q(q_out[5]) );
  DFFR_X1 \q_out_reg[4]  ( .D(N78), .CK(clock), .RN(n233), .Q(q_out[4]) );
  DFFR_X1 \q_out_reg[3]  ( .D(N77), .CK(clock), .RN(n233), .Q(q_out[3]) );
  DFFR_X1 \q_out_reg[2]  ( .D(N76), .CK(clock), .RN(n233), .Q(q_out[2]) );
  DFFR_X1 \q_out_reg[1]  ( .D(N75), .CK(clock), .RN(n233), .Q(q_out[1]) );
  DFFR_X1 \q_out_reg[0]  ( .D(n292), .CK(clock), .RN(n232), .Q(q_out[0]) );
  DFFR_X1 \result_reg[27]  ( .D(n312), .CK(clock), .RN(n232), .Q(result[27])
         );
  DFFR_X1 \result_reg[26]  ( .D(n311), .CK(clock), .RN(n232), .Q(result[26])
         );
  DFFR_X1 \result_reg[25]  ( .D(n310), .CK(clock), .RN(n232), .Q(result[25])
         );
  DFFR_X1 \result_reg[24]  ( .D(n309), .CK(clock), .RN(n232), .Q(result[24])
         );
  DFFR_X1 \result_reg[23]  ( .D(n308), .CK(clock), .RN(n232), .Q(result[23])
         );
  DFFR_X1 \result_reg[22]  ( .D(n307), .CK(clock), .RN(n232), .Q(result[22])
         );
  DFFR_X1 \result_reg[21]  ( .D(n306), .CK(clock), .RN(n232), .Q(result[21])
         );
  DFFR_X1 \result_reg[20]  ( .D(n305), .CK(clock), .RN(n232), .Q(result[20])
         );
  DFFR_X1 \result_reg[19]  ( .D(n304), .CK(clock), .RN(n232), .Q(result[19])
         );
  DFFR_X1 \result_reg[18]  ( .D(n303), .CK(clock), .RN(n232), .Q(result[18])
         );
  DFFR_X1 \result_reg[17]  ( .D(n302), .CK(clock), .RN(n232), .Q(result[17])
         );
  DFFR_X1 \result_reg[16]  ( .D(n301), .CK(clock), .RN(n231), .Q(result[16])
         );
  DFFR_X1 \result_reg[15]  ( .D(n300), .CK(clock), .RN(n231), .Q(result[15])
         );
  DFFR_X1 \result_reg[14]  ( .D(n299), .CK(clock), .RN(n231), .Q(result[14])
         );
  DFFR_X1 \result_reg[13]  ( .D(n298), .CK(clock), .RN(n231), .Q(result[13])
         );
  DFFR_X1 \result_reg[12]  ( .D(n297), .CK(clock), .RN(n231), .Q(result[12])
         );
  DFFR_X1 \result_reg[11]  ( .D(n296), .CK(clock), .RN(n231), .Q(result[11])
         );
  DFFR_X1 \result_reg[10]  ( .D(n295), .CK(clock), .RN(n231), .Q(result[10])
         );
  DFFR_X1 \result_reg[9]  ( .D(n294), .CK(clock), .RN(n231), .Q(result[9]) );
  DFFR_X1 \result_reg[8]  ( .D(n293), .CK(clock), .RN(n231), .Q(result[8]) );
  DFFR_X1 \result_reg[7]  ( .D(N53), .CK(clock), .RN(n231), .Q(result[7]) );
  DFFR_X1 \result_reg[6]  ( .D(N52), .CK(clock), .RN(n231), .Q(result[6]) );
  DFFR_X1 \result_reg[5]  ( .D(N51), .CK(clock), .RN(n231), .Q(result[5]) );
  DFFR_X1 \result_reg[4]  ( .D(N50), .CK(clock), .RN(n233), .Q(result[4]) );
  DFFR_X1 \result_reg[3]  ( .D(N49), .CK(clock), .RN(n230), .Q(result[3]) );
  DFFR_X1 \result_reg[2]  ( .D(N48), .CK(clock), .RN(n233), .Q(result[2]) );
  DFFR_X1 \result_reg[1]  ( .D(N47), .CK(clock), .RN(n233), .Q(result[1]) );
  DFFR_X1 \divisor_out_reg[19]  ( .D(N46), .CK(clock), .RN(n231), .Q(
        divisor_out[19]) );
  DFFR_X1 \divisor_out_reg[18]  ( .D(N45), .CK(clock), .RN(n230), .Q(
        divisor_out[18]) );
  DFFR_X1 \divisor_out_reg[17]  ( .D(N44), .CK(clock), .RN(n233), .Q(
        divisor_out[17]) );
  DFFR_X1 \divisor_out_reg[16]  ( .D(N43), .CK(clock), .RN(n232), .Q(
        divisor_out[16]) );
  DFFR_X1 \divisor_out_reg[15]  ( .D(N42), .CK(clock), .RN(n231), .Q(
        divisor_out[15]) );
  DFFR_X1 \divisor_out_reg[14]  ( .D(N41), .CK(clock), .RN(n230), .Q(
        divisor_out[14]) );
  DFFR_X1 \divisor_out_reg[13]  ( .D(N40), .CK(clock), .RN(n232), .Q(
        divisor_out[13]) );
  DFFR_X1 \divisor_out_reg[12]  ( .D(N39), .CK(clock), .RN(n233), .Q(
        divisor_out[12]) );
  DFFR_X1 \divisor_out_reg[11]  ( .D(N38), .CK(clock), .RN(n230), .Q(
        divisor_out[11]) );
  DFFR_X1 \divisor_out_reg[10]  ( .D(N37), .CK(clock), .RN(n230), .Q(
        divisor_out[10]) );
  DFFR_X1 \divisor_out_reg[9]  ( .D(N36), .CK(clock), .RN(n230), .Q(
        divisor_out[9]) );
  DFFR_X1 \divisor_out_reg[8]  ( .D(N35), .CK(clock), .RN(n230), .Q(
        divisor_out[8]) );
  DFFR_X1 \divisor_out_reg[7]  ( .D(N34), .CK(clock), .RN(n230), .Q(
        divisor_out[7]) );
  DFFR_X1 \divisor_out_reg[6]  ( .D(N33), .CK(clock), .RN(n230), .Q(
        divisor_out[6]) );
  DFFR_X1 \divisor_out_reg[5]  ( .D(N32), .CK(clock), .RN(n230), .Q(
        divisor_out[5]) );
  DFFR_X1 \divisor_out_reg[4]  ( .D(N31), .CK(clock), .RN(n230), .Q(
        divisor_out[4]) );
  DFFR_X1 \divisor_out_reg[3]  ( .D(N30), .CK(clock), .RN(n230), .Q(
        divisor_out[3]) );
  DFFR_X1 \divisor_out_reg[2]  ( .D(N29), .CK(clock), .RN(n230), .Q(
        divisor_out[2]) );
  DFFR_X1 \divisor_out_reg[1]  ( .D(N28), .CK(clock), .RN(n230), .Q(
        divisor_out[1]) );
  DFFR_X1 \divisor_out_reg[0]  ( .D(N27), .CK(clock), .RN(n230), .Q(
        divisor_out[0]) );
  AND2_X1 U47 ( .A1(start), .A2(q_in[6]), .ZN(N81) );
  AND2_X1 U48 ( .A1(q_in[5]), .A2(start), .ZN(N80) );
  AND2_X1 U49 ( .A1(q_in[4]), .A2(start), .ZN(N79) );
  AND2_X1 U50 ( .A1(q_in[3]), .A2(start), .ZN(N78) );
  AND2_X1 U51 ( .A1(q_in[2]), .A2(start), .ZN(N77) );
  AND2_X1 U52 ( .A1(q_in[1]), .A2(start), .ZN(N76) );
  AND2_X1 U53 ( .A1(q_in[0]), .A2(start), .ZN(N75) );
  AND2_X1 U56 ( .A1(divided[5]), .A2(start), .ZN(N52) );
  AND2_X1 U57 ( .A1(divided[4]), .A2(start), .ZN(N51) );
  AND2_X1 U58 ( .A1(divided[3]), .A2(start), .ZN(N50) );
  AND2_X1 U59 ( .A1(divided[2]), .A2(start), .ZN(N49) );
  AND2_X1 U60 ( .A1(divided[1]), .A2(start), .ZN(N48) );
  AND2_X1 U61 ( .A1(divided[0]), .A2(start), .ZN(N47) );
  AND2_X1 U62 ( .A1(divisor[19]), .A2(start), .ZN(N46) );
  AND2_X1 U63 ( .A1(divisor[18]), .A2(start), .ZN(N45) );
  AND2_X1 U64 ( .A1(divisor[17]), .A2(start), .ZN(N44) );
  AND2_X1 U65 ( .A1(divisor[16]), .A2(start), .ZN(N43) );
  AND2_X1 U66 ( .A1(divisor[15]), .A2(start), .ZN(N42) );
  AND2_X1 U67 ( .A1(divisor[14]), .A2(start), .ZN(N41) );
  AND2_X1 U68 ( .A1(divisor[13]), .A2(start), .ZN(N40) );
  divider_pipe_stage_6_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(result[0]) );
  INV_X4 U6 ( .A(n234), .ZN(n231) );
  INV_X4 U7 ( .A(n234), .ZN(n232) );
  INV_X4 U8 ( .A(n234), .ZN(n230) );
  INV_X4 U9 ( .A(n234), .ZN(n233) );
  INV_X4 U10 ( .A(reset_n), .ZN(n234) );
  NAND2_X2 U11 ( .A1(start), .A2(n235), .ZN(n276) );
  NAND2_X2 U12 ( .A1(start), .A2(n235), .ZN(n225) );
  NAND2_X2 U13 ( .A1(start), .A2(n235), .ZN(n226) );
  INV_X4 U14 ( .A(start), .ZN(n229) );
  NAND2_X2 U15 ( .A1(start), .A2(n236), .ZN(n227) );
  NAND2_X2 U16 ( .A1(start), .A2(n236), .ZN(n228) );
  XNOR2_X2 U17 ( .A(divided[27]), .B(stage_result[20]), .ZN(n236) );
  INV_X4 U18 ( .A(n236), .ZN(n235) );
  INV_X4 U19 ( .A(n276), .ZN(n292) );
  AND2_X1 U20 ( .A1(divided[6]), .A2(start), .ZN(N53) );
  NAND2_X2 U21 ( .A1(start), .A2(n236), .ZN(n278) );
  INV_X4 U22 ( .A(divided[7]), .ZN(n238) );
  INV_X4 U23 ( .A(stage_result[0]), .ZN(n237) );
  OAI22_X2 U24 ( .A1(n227), .A2(n238), .B1(n225), .B2(n237), .ZN(n293) );
  INV_X4 U25 ( .A(divided[8]), .ZN(n240) );
  INV_X4 U26 ( .A(stage_result[1]), .ZN(n239) );
  OAI22_X2 U27 ( .A1(n228), .A2(n240), .B1(n226), .B2(n239), .ZN(n294) );
  INV_X4 U28 ( .A(divided[9]), .ZN(n242) );
  INV_X4 U29 ( .A(stage_result[2]), .ZN(n241) );
  OAI22_X2 U30 ( .A1(n278), .A2(n242), .B1(n225), .B2(n241), .ZN(n295) );
  INV_X4 U31 ( .A(divided[10]), .ZN(n244) );
  INV_X4 U32 ( .A(stage_result[3]), .ZN(n243) );
  OAI22_X2 U33 ( .A1(n227), .A2(n244), .B1(n226), .B2(n243), .ZN(n296) );
  INV_X4 U34 ( .A(divided[11]), .ZN(n246) );
  INV_X4 U35 ( .A(stage_result[4]), .ZN(n245) );
  OAI22_X2 U36 ( .A1(n228), .A2(n246), .B1(n276), .B2(n245), .ZN(n297) );
  INV_X4 U37 ( .A(divided[12]), .ZN(n248) );
  INV_X4 U38 ( .A(stage_result[5]), .ZN(n247) );
  OAI22_X2 U39 ( .A1(n278), .A2(n248), .B1(n225), .B2(n247), .ZN(n298) );
  INV_X4 U40 ( .A(divided[13]), .ZN(n250) );
  INV_X4 U41 ( .A(stage_result[6]), .ZN(n249) );
  OAI22_X2 U42 ( .A1(n227), .A2(n250), .B1(n226), .B2(n249), .ZN(n299) );
  INV_X4 U43 ( .A(divided[14]), .ZN(n252) );
  INV_X4 U44 ( .A(stage_result[7]), .ZN(n251) );
  OAI22_X2 U45 ( .A1(n228), .A2(n252), .B1(n276), .B2(n251), .ZN(n300) );
  INV_X4 U46 ( .A(divided[15]), .ZN(n254) );
  INV_X4 U54 ( .A(stage_result[8]), .ZN(n253) );
  OAI22_X2 U55 ( .A1(n278), .A2(n254), .B1(n225), .B2(n253), .ZN(n301) );
  INV_X4 U69 ( .A(divided[16]), .ZN(n256) );
  INV_X4 U70 ( .A(stage_result[9]), .ZN(n255) );
  OAI22_X2 U71 ( .A1(n227), .A2(n256), .B1(n226), .B2(n255), .ZN(n302) );
  INV_X4 U72 ( .A(divided[17]), .ZN(n258) );
  INV_X4 U73 ( .A(stage_result[10]), .ZN(n257) );
  OAI22_X2 U74 ( .A1(n228), .A2(n258), .B1(n276), .B2(n257), .ZN(n303) );
  INV_X4 U75 ( .A(divided[18]), .ZN(n260) );
  INV_X4 U76 ( .A(stage_result[11]), .ZN(n259) );
  OAI22_X2 U77 ( .A1(n278), .A2(n260), .B1(n225), .B2(n259), .ZN(n304) );
  INV_X4 U78 ( .A(divided[19]), .ZN(n262) );
  INV_X4 U79 ( .A(stage_result[12]), .ZN(n261) );
  OAI22_X2 U80 ( .A1(n227), .A2(n262), .B1(n226), .B2(n261), .ZN(n305) );
  INV_X4 U81 ( .A(divided[20]), .ZN(n264) );
  INV_X4 U82 ( .A(stage_result[13]), .ZN(n263) );
  OAI22_X2 U83 ( .A1(n228), .A2(n264), .B1(n276), .B2(n263), .ZN(n306) );
  INV_X4 U84 ( .A(divided[21]), .ZN(n266) );
  INV_X4 U85 ( .A(stage_result[14]), .ZN(n265) );
  OAI22_X2 U86 ( .A1(n278), .A2(n266), .B1(n225), .B2(n265), .ZN(n307) );
  INV_X4 U87 ( .A(divided[22]), .ZN(n268) );
  INV_X4 U88 ( .A(stage_result[15]), .ZN(n267) );
  OAI22_X2 U89 ( .A1(n227), .A2(n268), .B1(n226), .B2(n267), .ZN(n308) );
  INV_X4 U90 ( .A(divided[23]), .ZN(n270) );
  INV_X4 U91 ( .A(stage_result[16]), .ZN(n269) );
  OAI22_X2 U92 ( .A1(n228), .A2(n270), .B1(n276), .B2(n269), .ZN(n309) );
  INV_X4 U93 ( .A(divided[24]), .ZN(n272) );
  INV_X4 U94 ( .A(stage_result[17]), .ZN(n271) );
  OAI22_X2 U95 ( .A1(n278), .A2(n272), .B1(n225), .B2(n271), .ZN(n310) );
  INV_X4 U96 ( .A(divided[25]), .ZN(n274) );
  INV_X4 U97 ( .A(stage_result[18]), .ZN(n273) );
  OAI22_X2 U98 ( .A1(n227), .A2(n274), .B1(n226), .B2(n273), .ZN(n311) );
  INV_X4 U99 ( .A(divided[26]), .ZN(n277) );
  INV_X4 U100 ( .A(stage_result[19]), .ZN(n275) );
  OAI22_X2 U101 ( .A1(n228), .A2(n277), .B1(n276), .B2(n275), .ZN(n312) );
  INV_X4 U102 ( .A(divisor[0]), .ZN(n279) );
  NOR2_X2 U103 ( .A1(n229), .A2(n279), .ZN(N27) );
  INV_X4 U104 ( .A(divisor[1]), .ZN(n280) );
  NOR2_X2 U105 ( .A1(n229), .A2(n280), .ZN(N28) );
  INV_X4 U106 ( .A(divisor[2]), .ZN(n281) );
  NOR2_X2 U107 ( .A1(n229), .A2(n281), .ZN(N29) );
  INV_X4 U108 ( .A(divisor[3]), .ZN(n282) );
  NOR2_X2 U109 ( .A1(n229), .A2(n282), .ZN(N30) );
  INV_X4 U110 ( .A(divisor[4]), .ZN(n283) );
  NOR2_X2 U111 ( .A1(n229), .A2(n283), .ZN(N31) );
  INV_X4 U112 ( .A(divisor[5]), .ZN(n284) );
  NOR2_X2 U113 ( .A1(n229), .A2(n284), .ZN(N32) );
  INV_X4 U114 ( .A(divisor[6]), .ZN(n285) );
  NOR2_X2 U115 ( .A1(n229), .A2(n285), .ZN(N33) );
  INV_X4 U116 ( .A(divisor[7]), .ZN(n286) );
  NOR2_X2 U117 ( .A1(n229), .A2(n286), .ZN(N34) );
  INV_X4 U118 ( .A(divisor[8]), .ZN(n287) );
  NOR2_X2 U119 ( .A1(n229), .A2(n287), .ZN(N35) );
  INV_X4 U120 ( .A(divisor[9]), .ZN(n288) );
  NOR2_X2 U121 ( .A1(n229), .A2(n288), .ZN(N36) );
  INV_X4 U122 ( .A(divisor[10]), .ZN(n289) );
  NOR2_X2 U123 ( .A1(n229), .A2(n289), .ZN(N37) );
  INV_X4 U124 ( .A(divisor[11]), .ZN(n290) );
  NOR2_X2 U125 ( .A1(n229), .A2(n290), .ZN(N38) );
  INV_X4 U126 ( .A(divisor[12]), .ZN(n291) );
  NOR2_X2 U127 ( .A1(n229), .A2(n291), .ZN(N39) );
endmodule


module divider_pipe_stage_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n110, n112, n114,
         n115, n116, n117, n118, n120, n121, n122;

  FA_X1 U2 ( .A(A[19]), .B(B[19]), .CI(n18), .CO(CO), .S(SUM[19]) );
  FA_X1 U3 ( .A(A[18]), .B(B[18]), .CI(n19), .CO(n18), .S(SUM[18]) );
  FA_X1 U4 ( .A(A[17]), .B(B[17]), .CI(n20), .CO(n19), .S(SUM[17]) );
  XOR2_X2 U5 ( .A(n1), .B(n23), .Z(SUM[16]) );
  NAND2_X2 U7 ( .A1(n107), .A2(n22), .ZN(n1) );
  NAND2_X2 U10 ( .A1(A[16]), .A2(B[16]), .ZN(n22) );
  XOR2_X2 U11 ( .A(n2), .B(n32), .Z(SUM[15]) );
  NAND2_X2 U15 ( .A1(n40), .A2(n28), .ZN(n26) );
  NAND2_X2 U19 ( .A1(n108), .A2(n31), .ZN(n2) );
  NAND2_X2 U22 ( .A1(A[15]), .A2(B[15]), .ZN(n31) );
  XNOR2_X2 U23 ( .A(n37), .B(n3), .ZN(SUM[14]) );
  NAND2_X2 U27 ( .A1(n33), .A2(n36), .ZN(n3) );
  NAND2_X2 U30 ( .A1(A[14]), .A2(B[14]), .ZN(n36) );
  XOR2_X2 U31 ( .A(n4), .B(n44), .Z(SUM[13]) );
  NAND2_X2 U37 ( .A1(n110), .A2(n43), .ZN(n4) );
  NAND2_X2 U40 ( .A1(A[13]), .A2(B[13]), .ZN(n43) );
  XOR2_X2 U41 ( .A(n5), .B(n49), .Z(SUM[12]) );
  NAND2_X2 U45 ( .A1(n45), .A2(n48), .ZN(n5) );
  NAND2_X2 U48 ( .A1(A[12]), .A2(B[12]), .ZN(n48) );
  XOR2_X2 U49 ( .A(n6), .B(n57), .Z(SUM[11]) );
  NAND2_X2 U52 ( .A1(n65), .A2(n53), .ZN(n51) );
  NAND2_X2 U56 ( .A1(n112), .A2(n56), .ZN(n6) );
  NAND2_X2 U59 ( .A1(A[11]), .A2(B[11]), .ZN(n56) );
  XNOR2_X2 U60 ( .A(n62), .B(n7), .ZN(SUM[10]) );
  NAND2_X2 U64 ( .A1(n58), .A2(n61), .ZN(n7) );
  NAND2_X2 U67 ( .A1(A[10]), .A2(B[10]), .ZN(n61) );
  XNOR2_X2 U68 ( .A(n69), .B(n8), .ZN(SUM[9]) );
  NAND2_X2 U74 ( .A1(n114), .A2(n68), .ZN(n8) );
  NAND2_X2 U77 ( .A1(A[9]), .A2(B[9]), .ZN(n68) );
  XOR2_X2 U78 ( .A(n9), .B(n72), .Z(SUM[8]) );
  NAND2_X2 U80 ( .A1(n115), .A2(n71), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[8]), .A2(B[8]), .ZN(n71) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[7]) );
  NAND2_X2 U87 ( .A1(n84), .A2(n76), .ZN(n74) );
  NAND2_X2 U91 ( .A1(n116), .A2(n79), .ZN(n10) );
  NAND2_X2 U94 ( .A1(A[7]), .A2(B[7]), .ZN(n79) );
  XOR2_X2 U95 ( .A(n11), .B(n83), .Z(SUM[6]) );
  NAND2_X2 U97 ( .A1(n117), .A2(n82), .ZN(n11) );
  NAND2_X2 U100 ( .A1(A[6]), .A2(B[6]), .ZN(n82) );
  XOR2_X2 U101 ( .A(n12), .B(n88), .Z(SUM[5]) );
  NAND2_X2 U105 ( .A1(n118), .A2(n87), .ZN(n12) );
  NAND2_X2 U108 ( .A1(A[5]), .A2(B[5]), .ZN(n87) );
  XNOR2_X2 U109 ( .A(n93), .B(n13), .ZN(SUM[4]) );
  NAND2_X2 U113 ( .A1(n89), .A2(n92), .ZN(n13) );
  NAND2_X2 U116 ( .A1(A[4]), .A2(B[4]), .ZN(n92) );
  XNOR2_X2 U117 ( .A(n99), .B(n14), .ZN(SUM[3]) );
  NAND2_X2 U122 ( .A1(n120), .A2(n98), .ZN(n14) );
  NAND2_X2 U125 ( .A1(A[3]), .A2(B[3]), .ZN(n98) );
  XOR2_X2 U126 ( .A(n15), .B(n102), .Z(SUM[2]) );
  NAND2_X2 U128 ( .A1(n121), .A2(n101), .ZN(n15) );
  NAND2_X2 U131 ( .A1(A[2]), .A2(B[2]), .ZN(n101) );
  XOR2_X2 U132 ( .A(n106), .B(n16), .Z(SUM[1]) );
  NAND2_X2 U135 ( .A1(n122), .A2(n105), .ZN(n16) );
  NAND2_X2 U138 ( .A1(A[1]), .A2(B[1]), .ZN(n105) );
  XNOR2_X2 U139 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U144 ( .B1(n73), .B2(n24), .A(n25), .ZN(n23) );
  NOR2_X2 U145 ( .A1(n51), .A2(n26), .ZN(n24) );
  OAI21_X2 U146 ( .B1(n52), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X2 U147 ( .B1(n49), .B2(n38), .A(n39), .ZN(n37) );
  OAI21_X2 U148 ( .B1(n72), .B2(n51), .A(n52), .ZN(n50) );
  AOI21_X2 U149 ( .B1(n93), .B2(n84), .A(n85), .ZN(n83) );
  OAI21_X2 U150 ( .B1(n72), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X2 U151 ( .B1(n53), .B2(n66), .A(n54), .ZN(n52) );
  OAI21_X2 U152 ( .B1(n55), .B2(n61), .A(n56), .ZN(n54) );
  AOI21_X2 U153 ( .B1(n95), .B2(n103), .A(n96), .ZN(n94) );
  NOR2_X2 U154 ( .A1(n100), .A2(n97), .ZN(n95) );
  OAI21_X2 U155 ( .B1(n97), .B2(n101), .A(n98), .ZN(n96) );
  OAI21_X2 U156 ( .B1(n86), .B2(n92), .A(n87), .ZN(n85) );
  OAI21_X2 U157 ( .B1(n94), .B2(n74), .A(n75), .ZN(n73) );
  AOI21_X2 U158 ( .B1(n76), .B2(n85), .A(n77), .ZN(n75) );
  NOR2_X2 U159 ( .A1(n81), .A2(n78), .ZN(n76) );
  AOI21_X2 U160 ( .B1(n28), .B2(n41), .A(n29), .ZN(n27) );
  OAI21_X2 U161 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  OAI21_X2 U162 ( .B1(n42), .B2(n48), .A(n43), .ZN(n41) );
  OAI21_X2 U163 ( .B1(n104), .B2(n106), .A(n105), .ZN(n103) );
  OAI21_X2 U164 ( .B1(n67), .B2(n71), .A(n68), .ZN(n66) );
  OAI21_X2 U165 ( .B1(n78), .B2(n82), .A(n79), .ZN(n77) );
  NOR2_X2 U166 ( .A1(n60), .A2(n55), .ZN(n53) );
  NOR2_X2 U167 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U168 ( .A1(n91), .A2(n86), .ZN(n84) );
  NOR2_X2 U169 ( .A1(n70), .A2(n67), .ZN(n65) );
  NOR2_X2 U170 ( .A1(n47), .A2(n42), .ZN(n40) );
  AOI21_X2 U171 ( .B1(n37), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U172 ( .B1(n93), .B2(n89), .A(n90), .ZN(n88) );
  AOI21_X2 U173 ( .B1(n62), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X2 U174 ( .B1(n50), .B2(n45), .A(n46), .ZN(n44) );
  OAI21_X2 U175 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X2 U176 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U177 ( .B1(n72), .B2(n70), .A(n71), .ZN(n69) );
  OAI21_X2 U178 ( .B1(n23), .B2(n21), .A(n22), .ZN(n20) );
  NOR2_X2 U179 ( .A1(A[3]), .A2(B[3]), .ZN(n97) );
  NOR2_X2 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n78) );
  NOR2_X2 U181 ( .A1(A[5]), .A2(B[5]), .ZN(n86) );
  NOR2_X2 U182 ( .A1(A[11]), .A2(B[11]), .ZN(n55) );
  NOR2_X2 U183 ( .A1(A[9]), .A2(B[9]), .ZN(n67) );
  NOR2_X2 U184 ( .A1(A[15]), .A2(B[15]), .ZN(n30) );
  NOR2_X2 U185 ( .A1(A[13]), .A2(B[13]), .ZN(n42) );
  NOR2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n100) );
  NOR2_X2 U187 ( .A1(A[6]), .A2(B[6]), .ZN(n81) );
  NOR2_X2 U188 ( .A1(A[8]), .A2(B[8]), .ZN(n70) );
  NOR2_X2 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n104) );
  NOR2_X2 U190 ( .A1(A[0]), .A2(B[0]), .ZN(n106) );
  NOR2_X2 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n91) );
  NOR2_X2 U192 ( .A1(A[10]), .A2(B[10]), .ZN(n60) );
  NOR2_X2 U193 ( .A1(A[12]), .A2(B[12]), .ZN(n47) );
  NOR2_X2 U194 ( .A1(A[14]), .A2(B[14]), .ZN(n35) );
  NOR2_X2 U195 ( .A1(A[16]), .A2(B[16]), .ZN(n21) );
  INV_X4 U196 ( .A(n94), .ZN(n93) );
  INV_X4 U197 ( .A(n92), .ZN(n90) );
  INV_X4 U198 ( .A(n73), .ZN(n72) );
  INV_X4 U199 ( .A(n66), .ZN(n64) );
  INV_X4 U200 ( .A(n65), .ZN(n63) );
  INV_X4 U201 ( .A(n61), .ZN(n59) );
  INV_X4 U202 ( .A(n50), .ZN(n49) );
  INV_X4 U203 ( .A(n48), .ZN(n46) );
  INV_X4 U204 ( .A(n41), .ZN(n39) );
  INV_X4 U205 ( .A(n40), .ZN(n38) );
  INV_X4 U206 ( .A(n36), .ZN(n34) );
  INV_X4 U207 ( .A(n104), .ZN(n122) );
  INV_X4 U208 ( .A(n100), .ZN(n121) );
  INV_X4 U209 ( .A(n97), .ZN(n120) );
  INV_X4 U210 ( .A(n91), .ZN(n89) );
  INV_X4 U211 ( .A(n86), .ZN(n118) );
  INV_X4 U212 ( .A(n81), .ZN(n117) );
  INV_X4 U213 ( .A(n78), .ZN(n116) );
  INV_X4 U214 ( .A(n70), .ZN(n115) );
  INV_X4 U215 ( .A(n67), .ZN(n114) );
  INV_X4 U216 ( .A(n60), .ZN(n58) );
  INV_X4 U217 ( .A(n55), .ZN(n112) );
  INV_X4 U218 ( .A(n47), .ZN(n45) );
  INV_X4 U219 ( .A(n42), .ZN(n110) );
  INV_X4 U220 ( .A(n35), .ZN(n33) );
  INV_X4 U221 ( .A(n30), .ZN(n108) );
  INV_X4 U222 ( .A(n21), .ZN(n107) );
  INV_X4 U223 ( .A(n103), .ZN(n102) );
endmodule


module divider_pipe_stage_5 ( clock, reset_n, start, divided, divisor, q_in, 
        start_out, divisor_out, result, q_out );
  input [27:0] divided;
  input [19:0] divisor;
  input [7:0] q_in;
  output [19:0] divisor_out;
  output [27:0] result;
  output [7:0] q_out;
  input clock, reset_n, start;
  output start_out;
  wire   N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N75,
         N76, N77, N78, N79, N80, N81, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313;
  wire   [20:0] stage_result;

  DFFR_X1 start_out_reg ( .D(n229), .CK(clock), .RN(n235), .Q(start_out) );
  DFFR_X1 \q_out_reg[7]  ( .D(N81), .CK(clock), .RN(n235), .Q(q_out[7]) );
  DFFR_X1 \q_out_reg[6]  ( .D(N80), .CK(clock), .RN(n235), .Q(q_out[6]) );
  DFFR_X1 \q_out_reg[5]  ( .D(N79), .CK(clock), .RN(n235), .Q(q_out[5]) );
  DFFR_X1 \q_out_reg[4]  ( .D(N78), .CK(clock), .RN(n235), .Q(q_out[4]) );
  DFFR_X1 \q_out_reg[3]  ( .D(N77), .CK(clock), .RN(n235), .Q(q_out[3]) );
  DFFR_X1 \q_out_reg[2]  ( .D(N76), .CK(clock), .RN(n235), .Q(q_out[2]) );
  DFFR_X1 \q_out_reg[1]  ( .D(N75), .CK(clock), .RN(n235), .Q(q_out[1]) );
  DFFR_X1 \q_out_reg[0]  ( .D(n293), .CK(clock), .RN(n234), .Q(q_out[0]) );
  DFFR_X1 \result_reg[27]  ( .D(n313), .CK(clock), .RN(n234), .Q(result[27])
         );
  DFFR_X1 \result_reg[26]  ( .D(n312), .CK(clock), .RN(n234), .Q(result[26])
         );
  DFFR_X1 \result_reg[25]  ( .D(n311), .CK(clock), .RN(n234), .Q(result[25])
         );
  DFFR_X1 \result_reg[24]  ( .D(n310), .CK(clock), .RN(n234), .Q(result[24])
         );
  DFFR_X1 \result_reg[23]  ( .D(n309), .CK(clock), .RN(n234), .Q(result[23])
         );
  DFFR_X1 \result_reg[22]  ( .D(n308), .CK(clock), .RN(n234), .Q(result[22])
         );
  DFFR_X1 \result_reg[21]  ( .D(n307), .CK(clock), .RN(n234), .Q(result[21])
         );
  DFFR_X1 \result_reg[20]  ( .D(n306), .CK(clock), .RN(n234), .Q(result[20])
         );
  DFFR_X1 \result_reg[19]  ( .D(n305), .CK(clock), .RN(n234), .Q(result[19])
         );
  DFFR_X1 \result_reg[18]  ( .D(n304), .CK(clock), .RN(n234), .Q(result[18])
         );
  DFFR_X1 \result_reg[17]  ( .D(n303), .CK(clock), .RN(n234), .Q(result[17])
         );
  DFFR_X1 \result_reg[16]  ( .D(n302), .CK(clock), .RN(reset_n), .Q(result[16]) );
  DFFR_X1 \result_reg[15]  ( .D(n301), .CK(clock), .RN(reset_n), .Q(result[15]) );
  DFFR_X1 \result_reg[14]  ( .D(n300), .CK(clock), .RN(n235), .Q(result[14])
         );
  DFFR_X1 \result_reg[13]  ( .D(n299), .CK(clock), .RN(reset_n), .Q(result[13]) );
  DFFR_X1 \result_reg[12]  ( .D(n298), .CK(clock), .RN(reset_n), .Q(result[12]) );
  DFFR_X1 \result_reg[11]  ( .D(n297), .CK(clock), .RN(reset_n), .Q(result[11]) );
  DFFR_X1 \result_reg[10]  ( .D(n296), .CK(clock), .RN(reset_n), .Q(result[10]) );
  DFFR_X1 \result_reg[9]  ( .D(n295), .CK(clock), .RN(n235), .Q(result[9]) );
  DFFR_X1 \result_reg[8]  ( .D(n294), .CK(clock), .RN(reset_n), .Q(result[8])
         );
  DFFR_X1 \result_reg[7]  ( .D(N53), .CK(clock), .RN(n234), .Q(result[7]) );
  DFFR_X1 \result_reg[6]  ( .D(N52), .CK(clock), .RN(n235), .Q(result[6]) );
  DFFR_X1 \result_reg[5]  ( .D(N51), .CK(clock), .RN(n235), .Q(result[5]) );
  DFFR_X1 \result_reg[4]  ( .D(N50), .CK(clock), .RN(n233), .Q(result[4]) );
  DFFR_X1 \result_reg[3]  ( .D(N49), .CK(clock), .RN(n233), .Q(result[3]) );
  DFFR_X1 \result_reg[2]  ( .D(N48), .CK(clock), .RN(n233), .Q(result[2]) );
  DFFR_X1 \result_reg[1]  ( .D(N47), .CK(clock), .RN(n233), .Q(result[1]) );
  DFFR_X1 \divisor_out_reg[19]  ( .D(N46), .CK(clock), .RN(n233), .Q(
        divisor_out[19]) );
  DFFR_X1 \divisor_out_reg[18]  ( .D(N45), .CK(clock), .RN(n233), .Q(
        divisor_out[18]) );
  DFFR_X1 \divisor_out_reg[17]  ( .D(N44), .CK(clock), .RN(n233), .Q(
        divisor_out[17]) );
  DFFR_X1 \divisor_out_reg[16]  ( .D(N43), .CK(clock), .RN(n233), .Q(
        divisor_out[16]) );
  DFFR_X1 \divisor_out_reg[15]  ( .D(N42), .CK(clock), .RN(n233), .Q(
        divisor_out[15]) );
  DFFR_X1 \divisor_out_reg[14]  ( .D(N41), .CK(clock), .RN(n233), .Q(
        divisor_out[14]) );
  DFFR_X1 \divisor_out_reg[13]  ( .D(N40), .CK(clock), .RN(n233), .Q(
        divisor_out[13]) );
  DFFR_X1 \divisor_out_reg[12]  ( .D(N39), .CK(clock), .RN(n233), .Q(
        divisor_out[12]) );
  DFFR_X1 \divisor_out_reg[11]  ( .D(N38), .CK(clock), .RN(n232), .Q(
        divisor_out[11]) );
  DFFR_X1 \divisor_out_reg[10]  ( .D(N37), .CK(clock), .RN(n232), .Q(
        divisor_out[10]) );
  DFFR_X1 \divisor_out_reg[9]  ( .D(N36), .CK(clock), .RN(n232), .Q(
        divisor_out[9]) );
  DFFR_X1 \divisor_out_reg[8]  ( .D(N35), .CK(clock), .RN(n232), .Q(
        divisor_out[8]) );
  DFFR_X1 \divisor_out_reg[7]  ( .D(N34), .CK(clock), .RN(n232), .Q(
        divisor_out[7]) );
  DFFR_X1 \divisor_out_reg[6]  ( .D(N33), .CK(clock), .RN(n232), .Q(
        divisor_out[6]) );
  DFFR_X1 \divisor_out_reg[5]  ( .D(N32), .CK(clock), .RN(n232), .Q(
        divisor_out[5]) );
  DFFR_X1 \divisor_out_reg[4]  ( .D(N31), .CK(clock), .RN(n232), .Q(
        divisor_out[4]) );
  DFFR_X1 \divisor_out_reg[3]  ( .D(N30), .CK(clock), .RN(n232), .Q(
        divisor_out[3]) );
  DFFR_X1 \divisor_out_reg[2]  ( .D(N29), .CK(clock), .RN(n232), .Q(
        divisor_out[2]) );
  DFFR_X1 \divisor_out_reg[1]  ( .D(N28), .CK(clock), .RN(n232), .Q(
        divisor_out[1]) );
  DFFR_X1 \divisor_out_reg[0]  ( .D(N27), .CK(clock), .RN(n232), .Q(
        divisor_out[0]) );
  AND2_X1 U47 ( .A1(n229), .A2(q_in[6]), .ZN(N81) );
  AND2_X1 U48 ( .A1(q_in[5]), .A2(n229), .ZN(N80) );
  AND2_X1 U49 ( .A1(q_in[4]), .A2(n229), .ZN(N79) );
  AND2_X1 U50 ( .A1(q_in[3]), .A2(n229), .ZN(N78) );
  AND2_X1 U51 ( .A1(q_in[2]), .A2(n229), .ZN(N77) );
  AND2_X1 U52 ( .A1(q_in[1]), .A2(n229), .ZN(N76) );
  AND2_X1 U53 ( .A1(q_in[0]), .A2(n229), .ZN(N75) );
  AND2_X1 U56 ( .A1(divided[5]), .A2(n229), .ZN(N52) );
  AND2_X1 U57 ( .A1(divided[4]), .A2(n229), .ZN(N51) );
  AND2_X1 U58 ( .A1(divided[3]), .A2(n229), .ZN(N50) );
  AND2_X1 U59 ( .A1(divided[2]), .A2(n229), .ZN(N49) );
  AND2_X1 U60 ( .A1(divided[1]), .A2(n229), .ZN(N48) );
  AND2_X1 U61 ( .A1(divided[0]), .A2(n229), .ZN(N47) );
  AND2_X1 U62 ( .A1(divisor[19]), .A2(n229), .ZN(N46) );
  AND2_X1 U63 ( .A1(divisor[18]), .A2(n229), .ZN(N45) );
  AND2_X1 U64 ( .A1(divisor[17]), .A2(n229), .ZN(N44) );
  AND2_X1 U65 ( .A1(divisor[16]), .A2(n229), .ZN(N43) );
  AND2_X1 U66 ( .A1(divisor[15]), .A2(n229), .ZN(N42) );
  AND2_X1 U67 ( .A1(divisor[14]), .A2(n229), .ZN(N41) );
  AND2_X1 U68 ( .A1(divisor[13]), .A2(n229), .ZN(N40) );
  divider_pipe_stage_5_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(result[0]) );
  INV_X4 U6 ( .A(n231), .ZN(n234) );
  INV_X4 U7 ( .A(n231), .ZN(n232) );
  INV_X4 U8 ( .A(n231), .ZN(n233) );
  INV_X4 U9 ( .A(n231), .ZN(n235) );
  INV_X4 U10 ( .A(reset_n), .ZN(n231) );
  NAND2_X2 U11 ( .A1(n229), .A2(n236), .ZN(n277) );
  NAND2_X2 U12 ( .A1(n229), .A2(n236), .ZN(n225) );
  NAND2_X2 U13 ( .A1(n229), .A2(n236), .ZN(n226) );
  INV_X4 U14 ( .A(n230), .ZN(n229) );
  INV_X4 U15 ( .A(start), .ZN(n230) );
  NAND2_X2 U16 ( .A1(n229), .A2(n237), .ZN(n227) );
  NAND2_X2 U17 ( .A1(n229), .A2(n237), .ZN(n228) );
  XNOR2_X2 U18 ( .A(divided[27]), .B(stage_result[20]), .ZN(n237) );
  INV_X4 U19 ( .A(n237), .ZN(n236) );
  INV_X4 U20 ( .A(n277), .ZN(n293) );
  AND2_X1 U21 ( .A1(divided[6]), .A2(n229), .ZN(N53) );
  NAND2_X2 U22 ( .A1(n229), .A2(n237), .ZN(n279) );
  INV_X4 U23 ( .A(divided[7]), .ZN(n239) );
  INV_X4 U24 ( .A(stage_result[0]), .ZN(n238) );
  OAI22_X2 U25 ( .A1(n227), .A2(n239), .B1(n225), .B2(n238), .ZN(n294) );
  INV_X4 U26 ( .A(divided[8]), .ZN(n241) );
  INV_X4 U27 ( .A(stage_result[1]), .ZN(n240) );
  OAI22_X2 U28 ( .A1(n228), .A2(n241), .B1(n226), .B2(n240), .ZN(n295) );
  INV_X4 U29 ( .A(divided[9]), .ZN(n243) );
  INV_X4 U30 ( .A(stage_result[2]), .ZN(n242) );
  OAI22_X2 U31 ( .A1(n279), .A2(n243), .B1(n225), .B2(n242), .ZN(n296) );
  INV_X4 U32 ( .A(divided[10]), .ZN(n245) );
  INV_X4 U33 ( .A(stage_result[3]), .ZN(n244) );
  OAI22_X2 U34 ( .A1(n227), .A2(n245), .B1(n226), .B2(n244), .ZN(n297) );
  INV_X4 U35 ( .A(divided[11]), .ZN(n247) );
  INV_X4 U36 ( .A(stage_result[4]), .ZN(n246) );
  OAI22_X2 U37 ( .A1(n228), .A2(n247), .B1(n277), .B2(n246), .ZN(n298) );
  INV_X4 U38 ( .A(divided[12]), .ZN(n249) );
  INV_X4 U39 ( .A(stage_result[5]), .ZN(n248) );
  OAI22_X2 U40 ( .A1(n279), .A2(n249), .B1(n225), .B2(n248), .ZN(n299) );
  INV_X4 U41 ( .A(divided[13]), .ZN(n251) );
  INV_X4 U42 ( .A(stage_result[6]), .ZN(n250) );
  OAI22_X2 U43 ( .A1(n227), .A2(n251), .B1(n226), .B2(n250), .ZN(n300) );
  INV_X4 U44 ( .A(divided[14]), .ZN(n253) );
  INV_X4 U45 ( .A(stage_result[7]), .ZN(n252) );
  OAI22_X2 U46 ( .A1(n228), .A2(n253), .B1(n277), .B2(n252), .ZN(n301) );
  INV_X4 U54 ( .A(divided[15]), .ZN(n255) );
  INV_X4 U55 ( .A(stage_result[8]), .ZN(n254) );
  OAI22_X2 U69 ( .A1(n279), .A2(n255), .B1(n225), .B2(n254), .ZN(n302) );
  INV_X4 U70 ( .A(divided[16]), .ZN(n257) );
  INV_X4 U71 ( .A(stage_result[9]), .ZN(n256) );
  OAI22_X2 U72 ( .A1(n227), .A2(n257), .B1(n226), .B2(n256), .ZN(n303) );
  INV_X4 U73 ( .A(divided[17]), .ZN(n259) );
  INV_X4 U74 ( .A(stage_result[10]), .ZN(n258) );
  OAI22_X2 U75 ( .A1(n228), .A2(n259), .B1(n277), .B2(n258), .ZN(n304) );
  INV_X4 U76 ( .A(divided[18]), .ZN(n261) );
  INV_X4 U77 ( .A(stage_result[11]), .ZN(n260) );
  OAI22_X2 U78 ( .A1(n279), .A2(n261), .B1(n225), .B2(n260), .ZN(n305) );
  INV_X4 U79 ( .A(divided[19]), .ZN(n263) );
  INV_X4 U80 ( .A(stage_result[12]), .ZN(n262) );
  OAI22_X2 U81 ( .A1(n227), .A2(n263), .B1(n226), .B2(n262), .ZN(n306) );
  INV_X4 U82 ( .A(divided[20]), .ZN(n265) );
  INV_X4 U83 ( .A(stage_result[13]), .ZN(n264) );
  OAI22_X2 U84 ( .A1(n228), .A2(n265), .B1(n277), .B2(n264), .ZN(n307) );
  INV_X4 U85 ( .A(divided[21]), .ZN(n267) );
  INV_X4 U86 ( .A(stage_result[14]), .ZN(n266) );
  OAI22_X2 U87 ( .A1(n279), .A2(n267), .B1(n225), .B2(n266), .ZN(n308) );
  INV_X4 U88 ( .A(divided[22]), .ZN(n269) );
  INV_X4 U89 ( .A(stage_result[15]), .ZN(n268) );
  OAI22_X2 U90 ( .A1(n227), .A2(n269), .B1(n226), .B2(n268), .ZN(n309) );
  INV_X4 U91 ( .A(divided[23]), .ZN(n271) );
  INV_X4 U92 ( .A(stage_result[16]), .ZN(n270) );
  OAI22_X2 U93 ( .A1(n228), .A2(n271), .B1(n277), .B2(n270), .ZN(n310) );
  INV_X4 U94 ( .A(divided[24]), .ZN(n273) );
  INV_X4 U95 ( .A(stage_result[17]), .ZN(n272) );
  OAI22_X2 U96 ( .A1(n279), .A2(n273), .B1(n225), .B2(n272), .ZN(n311) );
  INV_X4 U97 ( .A(divided[25]), .ZN(n275) );
  INV_X4 U98 ( .A(stage_result[18]), .ZN(n274) );
  OAI22_X2 U99 ( .A1(n227), .A2(n275), .B1(n226), .B2(n274), .ZN(n312) );
  INV_X4 U100 ( .A(divided[26]), .ZN(n278) );
  INV_X4 U101 ( .A(stage_result[19]), .ZN(n276) );
  OAI22_X2 U102 ( .A1(n228), .A2(n278), .B1(n277), .B2(n276), .ZN(n313) );
  INV_X4 U103 ( .A(divisor[0]), .ZN(n280) );
  NOR2_X2 U104 ( .A1(n230), .A2(n280), .ZN(N27) );
  INV_X4 U105 ( .A(divisor[1]), .ZN(n281) );
  NOR2_X2 U106 ( .A1(n230), .A2(n281), .ZN(N28) );
  INV_X4 U107 ( .A(divisor[2]), .ZN(n282) );
  NOR2_X2 U108 ( .A1(n230), .A2(n282), .ZN(N29) );
  INV_X4 U109 ( .A(divisor[3]), .ZN(n283) );
  NOR2_X2 U110 ( .A1(n230), .A2(n283), .ZN(N30) );
  INV_X4 U111 ( .A(divisor[4]), .ZN(n284) );
  NOR2_X2 U112 ( .A1(n230), .A2(n284), .ZN(N31) );
  INV_X4 U113 ( .A(divisor[5]), .ZN(n285) );
  NOR2_X2 U114 ( .A1(n230), .A2(n285), .ZN(N32) );
  INV_X4 U115 ( .A(divisor[6]), .ZN(n286) );
  NOR2_X2 U116 ( .A1(n230), .A2(n286), .ZN(N33) );
  INV_X4 U117 ( .A(divisor[7]), .ZN(n287) );
  NOR2_X2 U118 ( .A1(n230), .A2(n287), .ZN(N34) );
  INV_X4 U119 ( .A(divisor[8]), .ZN(n288) );
  NOR2_X2 U120 ( .A1(n230), .A2(n288), .ZN(N35) );
  INV_X4 U121 ( .A(divisor[9]), .ZN(n289) );
  NOR2_X2 U122 ( .A1(n230), .A2(n289), .ZN(N36) );
  INV_X4 U123 ( .A(divisor[10]), .ZN(n290) );
  NOR2_X2 U124 ( .A1(n230), .A2(n290), .ZN(N37) );
  INV_X4 U125 ( .A(divisor[11]), .ZN(n291) );
  NOR2_X2 U126 ( .A1(n230), .A2(n291), .ZN(N38) );
  INV_X4 U127 ( .A(divisor[12]), .ZN(n292) );
  NOR2_X2 U128 ( .A1(n230), .A2(n292), .ZN(N39) );
endmodule


module divider_pipe_stage_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n110, n112, n114,
         n115, n116, n117, n118, n120, n121, n122;

  FA_X1 U2 ( .A(A[19]), .B(B[19]), .CI(n18), .CO(CO), .S(SUM[19]) );
  FA_X1 U3 ( .A(A[18]), .B(B[18]), .CI(n19), .CO(n18), .S(SUM[18]) );
  FA_X1 U4 ( .A(A[17]), .B(B[17]), .CI(n20), .CO(n19), .S(SUM[17]) );
  XOR2_X2 U5 ( .A(n1), .B(n23), .Z(SUM[16]) );
  NAND2_X2 U7 ( .A1(n107), .A2(n22), .ZN(n1) );
  NAND2_X2 U10 ( .A1(A[16]), .A2(B[16]), .ZN(n22) );
  XOR2_X2 U11 ( .A(n2), .B(n32), .Z(SUM[15]) );
  NAND2_X2 U15 ( .A1(n40), .A2(n28), .ZN(n26) );
  NAND2_X2 U19 ( .A1(n108), .A2(n31), .ZN(n2) );
  NAND2_X2 U22 ( .A1(A[15]), .A2(B[15]), .ZN(n31) );
  XNOR2_X2 U23 ( .A(n37), .B(n3), .ZN(SUM[14]) );
  NAND2_X2 U27 ( .A1(n33), .A2(n36), .ZN(n3) );
  NAND2_X2 U30 ( .A1(A[14]), .A2(B[14]), .ZN(n36) );
  XOR2_X2 U31 ( .A(n4), .B(n44), .Z(SUM[13]) );
  NAND2_X2 U37 ( .A1(n110), .A2(n43), .ZN(n4) );
  NAND2_X2 U40 ( .A1(A[13]), .A2(B[13]), .ZN(n43) );
  XOR2_X2 U41 ( .A(n5), .B(n49), .Z(SUM[12]) );
  NAND2_X2 U45 ( .A1(n45), .A2(n48), .ZN(n5) );
  NAND2_X2 U48 ( .A1(A[12]), .A2(B[12]), .ZN(n48) );
  XOR2_X2 U49 ( .A(n6), .B(n57), .Z(SUM[11]) );
  NAND2_X2 U52 ( .A1(n65), .A2(n53), .ZN(n51) );
  NAND2_X2 U56 ( .A1(n112), .A2(n56), .ZN(n6) );
  NAND2_X2 U59 ( .A1(A[11]), .A2(B[11]), .ZN(n56) );
  XNOR2_X2 U60 ( .A(n62), .B(n7), .ZN(SUM[10]) );
  NAND2_X2 U64 ( .A1(n58), .A2(n61), .ZN(n7) );
  NAND2_X2 U67 ( .A1(A[10]), .A2(B[10]), .ZN(n61) );
  XNOR2_X2 U68 ( .A(n69), .B(n8), .ZN(SUM[9]) );
  NAND2_X2 U74 ( .A1(n114), .A2(n68), .ZN(n8) );
  NAND2_X2 U77 ( .A1(A[9]), .A2(B[9]), .ZN(n68) );
  XOR2_X2 U78 ( .A(n9), .B(n72), .Z(SUM[8]) );
  NAND2_X2 U80 ( .A1(n115), .A2(n71), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[8]), .A2(B[8]), .ZN(n71) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[7]) );
  NAND2_X2 U87 ( .A1(n84), .A2(n76), .ZN(n74) );
  NAND2_X2 U91 ( .A1(n116), .A2(n79), .ZN(n10) );
  NAND2_X2 U94 ( .A1(A[7]), .A2(B[7]), .ZN(n79) );
  XOR2_X2 U95 ( .A(n11), .B(n83), .Z(SUM[6]) );
  NAND2_X2 U97 ( .A1(n117), .A2(n82), .ZN(n11) );
  NAND2_X2 U100 ( .A1(A[6]), .A2(B[6]), .ZN(n82) );
  XOR2_X2 U101 ( .A(n12), .B(n88), .Z(SUM[5]) );
  NAND2_X2 U105 ( .A1(n118), .A2(n87), .ZN(n12) );
  NAND2_X2 U108 ( .A1(A[5]), .A2(B[5]), .ZN(n87) );
  XNOR2_X2 U109 ( .A(n93), .B(n13), .ZN(SUM[4]) );
  NAND2_X2 U113 ( .A1(n89), .A2(n92), .ZN(n13) );
  NAND2_X2 U116 ( .A1(A[4]), .A2(B[4]), .ZN(n92) );
  XNOR2_X2 U117 ( .A(n99), .B(n14), .ZN(SUM[3]) );
  NAND2_X2 U122 ( .A1(n120), .A2(n98), .ZN(n14) );
  NAND2_X2 U125 ( .A1(A[3]), .A2(B[3]), .ZN(n98) );
  XOR2_X2 U126 ( .A(n15), .B(n102), .Z(SUM[2]) );
  NAND2_X2 U128 ( .A1(n121), .A2(n101), .ZN(n15) );
  NAND2_X2 U131 ( .A1(A[2]), .A2(B[2]), .ZN(n101) );
  XOR2_X2 U132 ( .A(n106), .B(n16), .Z(SUM[1]) );
  NAND2_X2 U135 ( .A1(n122), .A2(n105), .ZN(n16) );
  NAND2_X2 U138 ( .A1(A[1]), .A2(B[1]), .ZN(n105) );
  XNOR2_X2 U139 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U144 ( .B1(n73), .B2(n24), .A(n25), .ZN(n23) );
  NOR2_X2 U145 ( .A1(n51), .A2(n26), .ZN(n24) );
  OAI21_X2 U146 ( .B1(n52), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X2 U147 ( .B1(n49), .B2(n38), .A(n39), .ZN(n37) );
  OAI21_X2 U148 ( .B1(n72), .B2(n51), .A(n52), .ZN(n50) );
  AOI21_X2 U149 ( .B1(n93), .B2(n84), .A(n85), .ZN(n83) );
  OAI21_X2 U150 ( .B1(n72), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X2 U151 ( .B1(n53), .B2(n66), .A(n54), .ZN(n52) );
  OAI21_X2 U152 ( .B1(n55), .B2(n61), .A(n56), .ZN(n54) );
  AOI21_X2 U153 ( .B1(n95), .B2(n103), .A(n96), .ZN(n94) );
  NOR2_X2 U154 ( .A1(n100), .A2(n97), .ZN(n95) );
  OAI21_X2 U155 ( .B1(n97), .B2(n101), .A(n98), .ZN(n96) );
  OAI21_X2 U156 ( .B1(n86), .B2(n92), .A(n87), .ZN(n85) );
  OAI21_X2 U157 ( .B1(n94), .B2(n74), .A(n75), .ZN(n73) );
  AOI21_X2 U158 ( .B1(n76), .B2(n85), .A(n77), .ZN(n75) );
  NOR2_X2 U159 ( .A1(n81), .A2(n78), .ZN(n76) );
  AOI21_X2 U160 ( .B1(n28), .B2(n41), .A(n29), .ZN(n27) );
  OAI21_X2 U161 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  OAI21_X2 U162 ( .B1(n42), .B2(n48), .A(n43), .ZN(n41) );
  OAI21_X2 U163 ( .B1(n104), .B2(n106), .A(n105), .ZN(n103) );
  OAI21_X2 U164 ( .B1(n67), .B2(n71), .A(n68), .ZN(n66) );
  OAI21_X2 U165 ( .B1(n78), .B2(n82), .A(n79), .ZN(n77) );
  NOR2_X2 U166 ( .A1(n60), .A2(n55), .ZN(n53) );
  NOR2_X2 U167 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U168 ( .A1(n91), .A2(n86), .ZN(n84) );
  NOR2_X2 U169 ( .A1(n70), .A2(n67), .ZN(n65) );
  NOR2_X2 U170 ( .A1(n47), .A2(n42), .ZN(n40) );
  AOI21_X2 U171 ( .B1(n37), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U172 ( .B1(n93), .B2(n89), .A(n90), .ZN(n88) );
  AOI21_X2 U173 ( .B1(n62), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X2 U174 ( .B1(n50), .B2(n45), .A(n46), .ZN(n44) );
  OAI21_X2 U175 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X2 U176 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U177 ( .B1(n72), .B2(n70), .A(n71), .ZN(n69) );
  OAI21_X2 U178 ( .B1(n23), .B2(n21), .A(n22), .ZN(n20) );
  NOR2_X2 U179 ( .A1(A[3]), .A2(B[3]), .ZN(n97) );
  NOR2_X2 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n78) );
  NOR2_X2 U181 ( .A1(A[5]), .A2(B[5]), .ZN(n86) );
  NOR2_X2 U182 ( .A1(A[11]), .A2(B[11]), .ZN(n55) );
  NOR2_X2 U183 ( .A1(A[9]), .A2(B[9]), .ZN(n67) );
  NOR2_X2 U184 ( .A1(A[15]), .A2(B[15]), .ZN(n30) );
  NOR2_X2 U185 ( .A1(A[13]), .A2(B[13]), .ZN(n42) );
  NOR2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n100) );
  NOR2_X2 U187 ( .A1(A[6]), .A2(B[6]), .ZN(n81) );
  NOR2_X2 U188 ( .A1(A[8]), .A2(B[8]), .ZN(n70) );
  NOR2_X2 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n104) );
  NOR2_X2 U190 ( .A1(A[0]), .A2(B[0]), .ZN(n106) );
  NOR2_X2 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n91) );
  NOR2_X2 U192 ( .A1(A[10]), .A2(B[10]), .ZN(n60) );
  NOR2_X2 U193 ( .A1(A[12]), .A2(B[12]), .ZN(n47) );
  NOR2_X2 U194 ( .A1(A[14]), .A2(B[14]), .ZN(n35) );
  NOR2_X2 U195 ( .A1(A[16]), .A2(B[16]), .ZN(n21) );
  INV_X4 U196 ( .A(n94), .ZN(n93) );
  INV_X4 U197 ( .A(n92), .ZN(n90) );
  INV_X4 U198 ( .A(n73), .ZN(n72) );
  INV_X4 U199 ( .A(n66), .ZN(n64) );
  INV_X4 U200 ( .A(n65), .ZN(n63) );
  INV_X4 U201 ( .A(n61), .ZN(n59) );
  INV_X4 U202 ( .A(n50), .ZN(n49) );
  INV_X4 U203 ( .A(n48), .ZN(n46) );
  INV_X4 U204 ( .A(n41), .ZN(n39) );
  INV_X4 U205 ( .A(n40), .ZN(n38) );
  INV_X4 U206 ( .A(n36), .ZN(n34) );
  INV_X4 U207 ( .A(n104), .ZN(n122) );
  INV_X4 U208 ( .A(n100), .ZN(n121) );
  INV_X4 U209 ( .A(n97), .ZN(n120) );
  INV_X4 U210 ( .A(n91), .ZN(n89) );
  INV_X4 U211 ( .A(n86), .ZN(n118) );
  INV_X4 U212 ( .A(n81), .ZN(n117) );
  INV_X4 U213 ( .A(n78), .ZN(n116) );
  INV_X4 U214 ( .A(n70), .ZN(n115) );
  INV_X4 U215 ( .A(n67), .ZN(n114) );
  INV_X4 U216 ( .A(n60), .ZN(n58) );
  INV_X4 U217 ( .A(n55), .ZN(n112) );
  INV_X4 U218 ( .A(n47), .ZN(n45) );
  INV_X4 U219 ( .A(n42), .ZN(n110) );
  INV_X4 U220 ( .A(n35), .ZN(n33) );
  INV_X4 U221 ( .A(n30), .ZN(n108) );
  INV_X4 U222 ( .A(n21), .ZN(n107) );
  INV_X4 U223 ( .A(n103), .ZN(n102) );
endmodule


module divider_pipe_stage_4 ( clock, reset_n, start, divided, divisor, q_in, 
        start_out, divisor_out, result, q_out );
  input [27:0] divided;
  input [19:0] divisor;
  input [7:0] q_in;
  output [19:0] divisor_out;
  output [27:0] result;
  output [7:0] q_out;
  input clock, reset_n, start;
  output start_out;
  wire   N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N75,
         N76, N77, N78, N79, N80, N81, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313;
  wire   [20:0] stage_result;

  DFFR_X1 start_out_reg ( .D(n229), .CK(clock), .RN(reset_n), .Q(start_out) );
  DFFR_X1 \q_out_reg[7]  ( .D(N81), .CK(clock), .RN(n231), .Q(q_out[7]) );
  DFFR_X1 \q_out_reg[6]  ( .D(N80), .CK(clock), .RN(n234), .Q(q_out[6]) );
  DFFR_X1 \q_out_reg[5]  ( .D(N79), .CK(clock), .RN(n233), .Q(q_out[5]) );
  DFFR_X1 \q_out_reg[4]  ( .D(N78), .CK(clock), .RN(n232), .Q(q_out[4]) );
  DFFR_X1 \q_out_reg[3]  ( .D(N77), .CK(clock), .RN(n231), .Q(q_out[3]) );
  DFFR_X1 \q_out_reg[2]  ( .D(N76), .CK(clock), .RN(n234), .Q(q_out[2]) );
  DFFR_X1 \q_out_reg[1]  ( .D(N75), .CK(clock), .RN(n233), .Q(q_out[1]) );
  DFFR_X1 \q_out_reg[0]  ( .D(n293), .CK(clock), .RN(n234), .Q(q_out[0]) );
  DFFR_X1 \result_reg[27]  ( .D(n313), .CK(clock), .RN(n234), .Q(result[27])
         );
  DFFR_X1 \result_reg[26]  ( .D(n312), .CK(clock), .RN(n234), .Q(result[26])
         );
  DFFR_X1 \result_reg[25]  ( .D(n311), .CK(clock), .RN(n234), .Q(result[25])
         );
  DFFR_X1 \result_reg[24]  ( .D(n310), .CK(clock), .RN(n234), .Q(result[24])
         );
  DFFR_X1 \result_reg[23]  ( .D(n309), .CK(clock), .RN(n234), .Q(result[23])
         );
  DFFR_X1 \result_reg[22]  ( .D(n308), .CK(clock), .RN(n234), .Q(result[22])
         );
  DFFR_X1 \result_reg[21]  ( .D(n307), .CK(clock), .RN(n234), .Q(result[21])
         );
  DFFR_X1 \result_reg[20]  ( .D(n306), .CK(clock), .RN(n234), .Q(result[20])
         );
  DFFR_X1 \result_reg[19]  ( .D(n305), .CK(clock), .RN(n234), .Q(result[19])
         );
  DFFR_X1 \result_reg[18]  ( .D(n304), .CK(clock), .RN(n234), .Q(result[18])
         );
  DFFR_X1 \result_reg[17]  ( .D(n303), .CK(clock), .RN(n234), .Q(result[17])
         );
  DFFR_X1 \result_reg[16]  ( .D(n302), .CK(clock), .RN(n233), .Q(result[16])
         );
  DFFR_X1 \result_reg[15]  ( .D(n301), .CK(clock), .RN(n233), .Q(result[15])
         );
  DFFR_X1 \result_reg[14]  ( .D(n300), .CK(clock), .RN(n233), .Q(result[14])
         );
  DFFR_X1 \result_reg[13]  ( .D(n299), .CK(clock), .RN(n233), .Q(result[13])
         );
  DFFR_X1 \result_reg[12]  ( .D(n298), .CK(clock), .RN(n233), .Q(result[12])
         );
  DFFR_X1 \result_reg[11]  ( .D(n297), .CK(clock), .RN(n233), .Q(result[11])
         );
  DFFR_X1 \result_reg[10]  ( .D(n296), .CK(clock), .RN(n233), .Q(result[10])
         );
  DFFR_X1 \result_reg[9]  ( .D(n295), .CK(clock), .RN(n233), .Q(result[9]) );
  DFFR_X1 \result_reg[8]  ( .D(n294), .CK(clock), .RN(n233), .Q(result[8]) );
  DFFR_X1 \result_reg[7]  ( .D(N53), .CK(clock), .RN(n233), .Q(result[7]) );
  DFFR_X1 \result_reg[6]  ( .D(N52), .CK(clock), .RN(n233), .Q(result[6]) );
  DFFR_X1 \result_reg[5]  ( .D(N51), .CK(clock), .RN(n233), .Q(result[5]) );
  DFFR_X1 \result_reg[4]  ( .D(N50), .CK(clock), .RN(n232), .Q(result[4]) );
  DFFR_X1 \result_reg[3]  ( .D(N49), .CK(clock), .RN(n232), .Q(result[3]) );
  DFFR_X1 \result_reg[2]  ( .D(N48), .CK(clock), .RN(n232), .Q(result[2]) );
  DFFR_X1 \result_reg[1]  ( .D(N47), .CK(clock), .RN(n232), .Q(result[1]) );
  DFFR_X1 \divisor_out_reg[19]  ( .D(N46), .CK(clock), .RN(n232), .Q(
        divisor_out[19]) );
  DFFR_X1 \divisor_out_reg[18]  ( .D(N45), .CK(clock), .RN(n232), .Q(
        divisor_out[18]) );
  DFFR_X1 \divisor_out_reg[17]  ( .D(N44), .CK(clock), .RN(n232), .Q(
        divisor_out[17]) );
  DFFR_X1 \divisor_out_reg[16]  ( .D(N43), .CK(clock), .RN(n232), .Q(
        divisor_out[16]) );
  DFFR_X1 \divisor_out_reg[15]  ( .D(N42), .CK(clock), .RN(n232), .Q(
        divisor_out[15]) );
  DFFR_X1 \divisor_out_reg[14]  ( .D(N41), .CK(clock), .RN(n232), .Q(
        divisor_out[14]) );
  DFFR_X1 \divisor_out_reg[13]  ( .D(N40), .CK(clock), .RN(n232), .Q(
        divisor_out[13]) );
  DFFR_X1 \divisor_out_reg[12]  ( .D(N39), .CK(clock), .RN(n232), .Q(
        divisor_out[12]) );
  DFFR_X1 \divisor_out_reg[11]  ( .D(N38), .CK(clock), .RN(n231), .Q(
        divisor_out[11]) );
  DFFR_X1 \divisor_out_reg[10]  ( .D(N37), .CK(clock), .RN(n231), .Q(
        divisor_out[10]) );
  DFFR_X1 \divisor_out_reg[9]  ( .D(N36), .CK(clock), .RN(n231), .Q(
        divisor_out[9]) );
  DFFR_X1 \divisor_out_reg[8]  ( .D(N35), .CK(clock), .RN(n231), .Q(
        divisor_out[8]) );
  DFFR_X1 \divisor_out_reg[7]  ( .D(N34), .CK(clock), .RN(n231), .Q(
        divisor_out[7]) );
  DFFR_X1 \divisor_out_reg[6]  ( .D(N33), .CK(clock), .RN(n231), .Q(
        divisor_out[6]) );
  DFFR_X1 \divisor_out_reg[5]  ( .D(N32), .CK(clock), .RN(n231), .Q(
        divisor_out[5]) );
  DFFR_X1 \divisor_out_reg[4]  ( .D(N31), .CK(clock), .RN(n231), .Q(
        divisor_out[4]) );
  DFFR_X1 \divisor_out_reg[3]  ( .D(N30), .CK(clock), .RN(n231), .Q(
        divisor_out[3]) );
  DFFR_X1 \divisor_out_reg[2]  ( .D(N29), .CK(clock), .RN(n231), .Q(
        divisor_out[2]) );
  DFFR_X1 \divisor_out_reg[1]  ( .D(N28), .CK(clock), .RN(n231), .Q(
        divisor_out[1]) );
  DFFR_X1 \divisor_out_reg[0]  ( .D(N27), .CK(clock), .RN(n231), .Q(
        divisor_out[0]) );
  AND2_X1 U47 ( .A1(n229), .A2(q_in[6]), .ZN(N81) );
  AND2_X1 U48 ( .A1(q_in[5]), .A2(n229), .ZN(N80) );
  AND2_X1 U49 ( .A1(q_in[4]), .A2(n229), .ZN(N79) );
  AND2_X1 U50 ( .A1(q_in[3]), .A2(n229), .ZN(N78) );
  AND2_X1 U51 ( .A1(q_in[2]), .A2(n229), .ZN(N77) );
  AND2_X1 U52 ( .A1(q_in[1]), .A2(n229), .ZN(N76) );
  AND2_X1 U53 ( .A1(q_in[0]), .A2(n229), .ZN(N75) );
  AND2_X1 U56 ( .A1(divided[5]), .A2(n229), .ZN(N52) );
  AND2_X1 U57 ( .A1(divided[4]), .A2(n229), .ZN(N51) );
  AND2_X1 U58 ( .A1(divided[3]), .A2(n229), .ZN(N50) );
  AND2_X1 U59 ( .A1(divided[2]), .A2(n229), .ZN(N49) );
  AND2_X1 U60 ( .A1(divided[1]), .A2(n229), .ZN(N48) );
  AND2_X1 U61 ( .A1(divided[0]), .A2(n229), .ZN(N47) );
  AND2_X1 U62 ( .A1(divisor[19]), .A2(n229), .ZN(N46) );
  AND2_X1 U63 ( .A1(divisor[18]), .A2(n229), .ZN(N45) );
  AND2_X1 U64 ( .A1(divisor[17]), .A2(n229), .ZN(N44) );
  AND2_X1 U65 ( .A1(divisor[16]), .A2(n229), .ZN(N43) );
  AND2_X1 U66 ( .A1(divisor[15]), .A2(n229), .ZN(N42) );
  AND2_X1 U67 ( .A1(divisor[14]), .A2(n229), .ZN(N41) );
  AND2_X1 U68 ( .A1(divisor[13]), .A2(n229), .ZN(N40) );
  divider_pipe_stage_4_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(result[0]) );
  INV_X4 U6 ( .A(n235), .ZN(n233) );
  INV_X4 U7 ( .A(n235), .ZN(n234) );
  INV_X4 U8 ( .A(n235), .ZN(n231) );
  INV_X4 U9 ( .A(n235), .ZN(n232) );
  INV_X4 U10 ( .A(reset_n), .ZN(n235) );
  NAND2_X2 U11 ( .A1(n229), .A2(n236), .ZN(n277) );
  NAND2_X2 U12 ( .A1(n229), .A2(n236), .ZN(n225) );
  NAND2_X2 U13 ( .A1(n229), .A2(n236), .ZN(n226) );
  INV_X4 U14 ( .A(n230), .ZN(n229) );
  INV_X4 U15 ( .A(start), .ZN(n230) );
  NAND2_X2 U16 ( .A1(n229), .A2(n237), .ZN(n227) );
  NAND2_X2 U17 ( .A1(n229), .A2(n237), .ZN(n228) );
  XNOR2_X2 U18 ( .A(divided[27]), .B(stage_result[20]), .ZN(n237) );
  INV_X4 U19 ( .A(n237), .ZN(n236) );
  INV_X4 U20 ( .A(n277), .ZN(n293) );
  AND2_X1 U21 ( .A1(divided[6]), .A2(n229), .ZN(N53) );
  NAND2_X2 U22 ( .A1(n229), .A2(n237), .ZN(n279) );
  INV_X4 U23 ( .A(divided[7]), .ZN(n239) );
  INV_X4 U24 ( .A(stage_result[0]), .ZN(n238) );
  OAI22_X2 U25 ( .A1(n227), .A2(n239), .B1(n225), .B2(n238), .ZN(n294) );
  INV_X4 U26 ( .A(divided[8]), .ZN(n241) );
  INV_X4 U27 ( .A(stage_result[1]), .ZN(n240) );
  OAI22_X2 U28 ( .A1(n228), .A2(n241), .B1(n226), .B2(n240), .ZN(n295) );
  INV_X4 U29 ( .A(divided[9]), .ZN(n243) );
  INV_X4 U30 ( .A(stage_result[2]), .ZN(n242) );
  OAI22_X2 U31 ( .A1(n279), .A2(n243), .B1(n225), .B2(n242), .ZN(n296) );
  INV_X4 U32 ( .A(divided[10]), .ZN(n245) );
  INV_X4 U33 ( .A(stage_result[3]), .ZN(n244) );
  OAI22_X2 U34 ( .A1(n227), .A2(n245), .B1(n226), .B2(n244), .ZN(n297) );
  INV_X4 U35 ( .A(divided[11]), .ZN(n247) );
  INV_X4 U36 ( .A(stage_result[4]), .ZN(n246) );
  OAI22_X2 U37 ( .A1(n228), .A2(n247), .B1(n277), .B2(n246), .ZN(n298) );
  INV_X4 U38 ( .A(divided[12]), .ZN(n249) );
  INV_X4 U39 ( .A(stage_result[5]), .ZN(n248) );
  OAI22_X2 U40 ( .A1(n279), .A2(n249), .B1(n225), .B2(n248), .ZN(n299) );
  INV_X4 U41 ( .A(divided[13]), .ZN(n251) );
  INV_X4 U42 ( .A(stage_result[6]), .ZN(n250) );
  OAI22_X2 U43 ( .A1(n227), .A2(n251), .B1(n226), .B2(n250), .ZN(n300) );
  INV_X4 U44 ( .A(divided[14]), .ZN(n253) );
  INV_X4 U45 ( .A(stage_result[7]), .ZN(n252) );
  OAI22_X2 U46 ( .A1(n228), .A2(n253), .B1(n277), .B2(n252), .ZN(n301) );
  INV_X4 U54 ( .A(divided[15]), .ZN(n255) );
  INV_X4 U55 ( .A(stage_result[8]), .ZN(n254) );
  OAI22_X2 U69 ( .A1(n279), .A2(n255), .B1(n225), .B2(n254), .ZN(n302) );
  INV_X4 U70 ( .A(divided[16]), .ZN(n257) );
  INV_X4 U71 ( .A(stage_result[9]), .ZN(n256) );
  OAI22_X2 U72 ( .A1(n227), .A2(n257), .B1(n226), .B2(n256), .ZN(n303) );
  INV_X4 U73 ( .A(divided[17]), .ZN(n259) );
  INV_X4 U74 ( .A(stage_result[10]), .ZN(n258) );
  OAI22_X2 U75 ( .A1(n228), .A2(n259), .B1(n277), .B2(n258), .ZN(n304) );
  INV_X4 U76 ( .A(divided[18]), .ZN(n261) );
  INV_X4 U77 ( .A(stage_result[11]), .ZN(n260) );
  OAI22_X2 U78 ( .A1(n279), .A2(n261), .B1(n225), .B2(n260), .ZN(n305) );
  INV_X4 U79 ( .A(divided[19]), .ZN(n263) );
  INV_X4 U80 ( .A(stage_result[12]), .ZN(n262) );
  OAI22_X2 U81 ( .A1(n227), .A2(n263), .B1(n226), .B2(n262), .ZN(n306) );
  INV_X4 U82 ( .A(divided[20]), .ZN(n265) );
  INV_X4 U83 ( .A(stage_result[13]), .ZN(n264) );
  OAI22_X2 U84 ( .A1(n228), .A2(n265), .B1(n277), .B2(n264), .ZN(n307) );
  INV_X4 U85 ( .A(divided[21]), .ZN(n267) );
  INV_X4 U86 ( .A(stage_result[14]), .ZN(n266) );
  OAI22_X2 U87 ( .A1(n279), .A2(n267), .B1(n225), .B2(n266), .ZN(n308) );
  INV_X4 U88 ( .A(divided[22]), .ZN(n269) );
  INV_X4 U89 ( .A(stage_result[15]), .ZN(n268) );
  OAI22_X2 U90 ( .A1(n227), .A2(n269), .B1(n226), .B2(n268), .ZN(n309) );
  INV_X4 U91 ( .A(divided[23]), .ZN(n271) );
  INV_X4 U92 ( .A(stage_result[16]), .ZN(n270) );
  OAI22_X2 U93 ( .A1(n228), .A2(n271), .B1(n277), .B2(n270), .ZN(n310) );
  INV_X4 U94 ( .A(divided[24]), .ZN(n273) );
  INV_X4 U95 ( .A(stage_result[17]), .ZN(n272) );
  OAI22_X2 U96 ( .A1(n279), .A2(n273), .B1(n225), .B2(n272), .ZN(n311) );
  INV_X4 U97 ( .A(divided[25]), .ZN(n275) );
  INV_X4 U98 ( .A(stage_result[18]), .ZN(n274) );
  OAI22_X2 U99 ( .A1(n227), .A2(n275), .B1(n226), .B2(n274), .ZN(n312) );
  INV_X4 U100 ( .A(divided[26]), .ZN(n278) );
  INV_X4 U101 ( .A(stage_result[19]), .ZN(n276) );
  OAI22_X2 U102 ( .A1(n228), .A2(n278), .B1(n277), .B2(n276), .ZN(n313) );
  INV_X4 U103 ( .A(divisor[0]), .ZN(n280) );
  NOR2_X2 U104 ( .A1(n230), .A2(n280), .ZN(N27) );
  INV_X4 U105 ( .A(divisor[1]), .ZN(n281) );
  NOR2_X2 U106 ( .A1(n230), .A2(n281), .ZN(N28) );
  INV_X4 U107 ( .A(divisor[2]), .ZN(n282) );
  NOR2_X2 U108 ( .A1(n230), .A2(n282), .ZN(N29) );
  INV_X4 U109 ( .A(divisor[3]), .ZN(n283) );
  NOR2_X2 U110 ( .A1(n230), .A2(n283), .ZN(N30) );
  INV_X4 U111 ( .A(divisor[4]), .ZN(n284) );
  NOR2_X2 U112 ( .A1(n230), .A2(n284), .ZN(N31) );
  INV_X4 U113 ( .A(divisor[5]), .ZN(n285) );
  NOR2_X2 U114 ( .A1(n230), .A2(n285), .ZN(N32) );
  INV_X4 U115 ( .A(divisor[6]), .ZN(n286) );
  NOR2_X2 U116 ( .A1(n230), .A2(n286), .ZN(N33) );
  INV_X4 U117 ( .A(divisor[7]), .ZN(n287) );
  NOR2_X2 U118 ( .A1(n230), .A2(n287), .ZN(N34) );
  INV_X4 U119 ( .A(divisor[8]), .ZN(n288) );
  NOR2_X2 U120 ( .A1(n230), .A2(n288), .ZN(N35) );
  INV_X4 U121 ( .A(divisor[9]), .ZN(n289) );
  NOR2_X2 U122 ( .A1(n230), .A2(n289), .ZN(N36) );
  INV_X4 U123 ( .A(divisor[10]), .ZN(n290) );
  NOR2_X2 U124 ( .A1(n230), .A2(n290), .ZN(N37) );
  INV_X4 U125 ( .A(divisor[11]), .ZN(n291) );
  NOR2_X2 U126 ( .A1(n230), .A2(n291), .ZN(N38) );
  INV_X4 U127 ( .A(divisor[12]), .ZN(n292) );
  NOR2_X2 U128 ( .A1(n230), .A2(n292), .ZN(N39) );
endmodule


module divider_pipe_stage_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n110, n112, n114,
         n115, n116, n117, n118, n120, n121, n122;

  FA_X1 U2 ( .A(A[19]), .B(B[19]), .CI(n18), .CO(CO), .S(SUM[19]) );
  FA_X1 U3 ( .A(A[18]), .B(B[18]), .CI(n19), .CO(n18), .S(SUM[18]) );
  FA_X1 U4 ( .A(A[17]), .B(B[17]), .CI(n20), .CO(n19), .S(SUM[17]) );
  XOR2_X2 U5 ( .A(n1), .B(n23), .Z(SUM[16]) );
  NAND2_X2 U7 ( .A1(n107), .A2(n22), .ZN(n1) );
  NAND2_X2 U10 ( .A1(A[16]), .A2(B[16]), .ZN(n22) );
  XOR2_X2 U11 ( .A(n2), .B(n32), .Z(SUM[15]) );
  NAND2_X2 U15 ( .A1(n40), .A2(n28), .ZN(n26) );
  NAND2_X2 U19 ( .A1(n108), .A2(n31), .ZN(n2) );
  NAND2_X2 U22 ( .A1(A[15]), .A2(B[15]), .ZN(n31) );
  XNOR2_X2 U23 ( .A(n37), .B(n3), .ZN(SUM[14]) );
  NAND2_X2 U27 ( .A1(n33), .A2(n36), .ZN(n3) );
  NAND2_X2 U30 ( .A1(A[14]), .A2(B[14]), .ZN(n36) );
  XOR2_X2 U31 ( .A(n4), .B(n44), .Z(SUM[13]) );
  NAND2_X2 U37 ( .A1(n110), .A2(n43), .ZN(n4) );
  NAND2_X2 U40 ( .A1(A[13]), .A2(B[13]), .ZN(n43) );
  XOR2_X2 U41 ( .A(n5), .B(n49), .Z(SUM[12]) );
  NAND2_X2 U45 ( .A1(n45), .A2(n48), .ZN(n5) );
  NAND2_X2 U48 ( .A1(A[12]), .A2(B[12]), .ZN(n48) );
  XOR2_X2 U49 ( .A(n6), .B(n57), .Z(SUM[11]) );
  NAND2_X2 U52 ( .A1(n65), .A2(n53), .ZN(n51) );
  NAND2_X2 U56 ( .A1(n112), .A2(n56), .ZN(n6) );
  NAND2_X2 U59 ( .A1(A[11]), .A2(B[11]), .ZN(n56) );
  XNOR2_X2 U60 ( .A(n62), .B(n7), .ZN(SUM[10]) );
  NAND2_X2 U64 ( .A1(n58), .A2(n61), .ZN(n7) );
  NAND2_X2 U67 ( .A1(A[10]), .A2(B[10]), .ZN(n61) );
  XNOR2_X2 U68 ( .A(n69), .B(n8), .ZN(SUM[9]) );
  NAND2_X2 U74 ( .A1(n114), .A2(n68), .ZN(n8) );
  NAND2_X2 U77 ( .A1(A[9]), .A2(B[9]), .ZN(n68) );
  XOR2_X2 U78 ( .A(n9), .B(n72), .Z(SUM[8]) );
  NAND2_X2 U80 ( .A1(n115), .A2(n71), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[8]), .A2(B[8]), .ZN(n71) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[7]) );
  NAND2_X2 U87 ( .A1(n84), .A2(n76), .ZN(n74) );
  NAND2_X2 U91 ( .A1(n116), .A2(n79), .ZN(n10) );
  NAND2_X2 U94 ( .A1(A[7]), .A2(B[7]), .ZN(n79) );
  XOR2_X2 U95 ( .A(n11), .B(n83), .Z(SUM[6]) );
  NAND2_X2 U97 ( .A1(n117), .A2(n82), .ZN(n11) );
  NAND2_X2 U100 ( .A1(A[6]), .A2(B[6]), .ZN(n82) );
  XOR2_X2 U101 ( .A(n12), .B(n88), .Z(SUM[5]) );
  NAND2_X2 U105 ( .A1(n118), .A2(n87), .ZN(n12) );
  NAND2_X2 U108 ( .A1(A[5]), .A2(B[5]), .ZN(n87) );
  XNOR2_X2 U109 ( .A(n93), .B(n13), .ZN(SUM[4]) );
  NAND2_X2 U113 ( .A1(n89), .A2(n92), .ZN(n13) );
  NAND2_X2 U116 ( .A1(A[4]), .A2(B[4]), .ZN(n92) );
  XNOR2_X2 U117 ( .A(n99), .B(n14), .ZN(SUM[3]) );
  NAND2_X2 U122 ( .A1(n120), .A2(n98), .ZN(n14) );
  NAND2_X2 U125 ( .A1(A[3]), .A2(B[3]), .ZN(n98) );
  XOR2_X2 U126 ( .A(n15), .B(n102), .Z(SUM[2]) );
  NAND2_X2 U128 ( .A1(n121), .A2(n101), .ZN(n15) );
  NAND2_X2 U131 ( .A1(A[2]), .A2(B[2]), .ZN(n101) );
  XOR2_X2 U132 ( .A(n106), .B(n16), .Z(SUM[1]) );
  NAND2_X2 U135 ( .A1(n122), .A2(n105), .ZN(n16) );
  NAND2_X2 U138 ( .A1(A[1]), .A2(B[1]), .ZN(n105) );
  XNOR2_X2 U139 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U144 ( .B1(n73), .B2(n24), .A(n25), .ZN(n23) );
  NOR2_X2 U145 ( .A1(n51), .A2(n26), .ZN(n24) );
  OAI21_X2 U146 ( .B1(n52), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X2 U147 ( .B1(n49), .B2(n38), .A(n39), .ZN(n37) );
  OAI21_X2 U148 ( .B1(n72), .B2(n51), .A(n52), .ZN(n50) );
  AOI21_X2 U149 ( .B1(n93), .B2(n84), .A(n85), .ZN(n83) );
  OAI21_X2 U150 ( .B1(n72), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X2 U151 ( .B1(n53), .B2(n66), .A(n54), .ZN(n52) );
  OAI21_X2 U152 ( .B1(n55), .B2(n61), .A(n56), .ZN(n54) );
  AOI21_X2 U153 ( .B1(n95), .B2(n103), .A(n96), .ZN(n94) );
  NOR2_X2 U154 ( .A1(n100), .A2(n97), .ZN(n95) );
  OAI21_X2 U155 ( .B1(n97), .B2(n101), .A(n98), .ZN(n96) );
  OAI21_X2 U156 ( .B1(n86), .B2(n92), .A(n87), .ZN(n85) );
  OAI21_X2 U157 ( .B1(n94), .B2(n74), .A(n75), .ZN(n73) );
  AOI21_X2 U158 ( .B1(n76), .B2(n85), .A(n77), .ZN(n75) );
  NOR2_X2 U159 ( .A1(n81), .A2(n78), .ZN(n76) );
  AOI21_X2 U160 ( .B1(n28), .B2(n41), .A(n29), .ZN(n27) );
  OAI21_X2 U161 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  OAI21_X2 U162 ( .B1(n42), .B2(n48), .A(n43), .ZN(n41) );
  OAI21_X2 U163 ( .B1(n104), .B2(n106), .A(n105), .ZN(n103) );
  OAI21_X2 U164 ( .B1(n67), .B2(n71), .A(n68), .ZN(n66) );
  OAI21_X2 U165 ( .B1(n78), .B2(n82), .A(n79), .ZN(n77) );
  NOR2_X2 U166 ( .A1(n60), .A2(n55), .ZN(n53) );
  NOR2_X2 U167 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U168 ( .A1(n91), .A2(n86), .ZN(n84) );
  NOR2_X2 U169 ( .A1(n70), .A2(n67), .ZN(n65) );
  NOR2_X2 U170 ( .A1(n47), .A2(n42), .ZN(n40) );
  AOI21_X2 U171 ( .B1(n37), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U172 ( .B1(n93), .B2(n89), .A(n90), .ZN(n88) );
  AOI21_X2 U173 ( .B1(n62), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X2 U174 ( .B1(n50), .B2(n45), .A(n46), .ZN(n44) );
  OAI21_X2 U175 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X2 U176 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U177 ( .B1(n72), .B2(n70), .A(n71), .ZN(n69) );
  OAI21_X2 U178 ( .B1(n23), .B2(n21), .A(n22), .ZN(n20) );
  NOR2_X2 U179 ( .A1(A[3]), .A2(B[3]), .ZN(n97) );
  NOR2_X2 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n78) );
  NOR2_X2 U181 ( .A1(A[5]), .A2(B[5]), .ZN(n86) );
  NOR2_X2 U182 ( .A1(A[11]), .A2(B[11]), .ZN(n55) );
  NOR2_X2 U183 ( .A1(A[9]), .A2(B[9]), .ZN(n67) );
  NOR2_X2 U184 ( .A1(A[15]), .A2(B[15]), .ZN(n30) );
  NOR2_X2 U185 ( .A1(A[13]), .A2(B[13]), .ZN(n42) );
  NOR2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n100) );
  NOR2_X2 U187 ( .A1(A[6]), .A2(B[6]), .ZN(n81) );
  NOR2_X2 U188 ( .A1(A[8]), .A2(B[8]), .ZN(n70) );
  NOR2_X2 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n104) );
  NOR2_X2 U190 ( .A1(A[0]), .A2(B[0]), .ZN(n106) );
  NOR2_X2 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n91) );
  NOR2_X2 U192 ( .A1(A[10]), .A2(B[10]), .ZN(n60) );
  NOR2_X2 U193 ( .A1(A[12]), .A2(B[12]), .ZN(n47) );
  NOR2_X2 U194 ( .A1(A[14]), .A2(B[14]), .ZN(n35) );
  NOR2_X2 U195 ( .A1(A[16]), .A2(B[16]), .ZN(n21) );
  INV_X4 U196 ( .A(n94), .ZN(n93) );
  INV_X4 U197 ( .A(n92), .ZN(n90) );
  INV_X4 U198 ( .A(n73), .ZN(n72) );
  INV_X4 U199 ( .A(n66), .ZN(n64) );
  INV_X4 U200 ( .A(n65), .ZN(n63) );
  INV_X4 U201 ( .A(n61), .ZN(n59) );
  INV_X4 U202 ( .A(n50), .ZN(n49) );
  INV_X4 U203 ( .A(n48), .ZN(n46) );
  INV_X4 U204 ( .A(n41), .ZN(n39) );
  INV_X4 U205 ( .A(n40), .ZN(n38) );
  INV_X4 U206 ( .A(n36), .ZN(n34) );
  INV_X4 U207 ( .A(n104), .ZN(n122) );
  INV_X4 U208 ( .A(n100), .ZN(n121) );
  INV_X4 U209 ( .A(n97), .ZN(n120) );
  INV_X4 U210 ( .A(n91), .ZN(n89) );
  INV_X4 U211 ( .A(n86), .ZN(n118) );
  INV_X4 U212 ( .A(n81), .ZN(n117) );
  INV_X4 U213 ( .A(n78), .ZN(n116) );
  INV_X4 U214 ( .A(n70), .ZN(n115) );
  INV_X4 U215 ( .A(n67), .ZN(n114) );
  INV_X4 U216 ( .A(n60), .ZN(n58) );
  INV_X4 U217 ( .A(n55), .ZN(n112) );
  INV_X4 U218 ( .A(n47), .ZN(n45) );
  INV_X4 U219 ( .A(n42), .ZN(n110) );
  INV_X4 U220 ( .A(n35), .ZN(n33) );
  INV_X4 U221 ( .A(n30), .ZN(n108) );
  INV_X4 U222 ( .A(n21), .ZN(n107) );
  INV_X4 U223 ( .A(n103), .ZN(n102) );
endmodule


module divider_pipe_stage_3 ( clock, reset_n, start, divided, divisor, q_in, 
        start_out, divisor_out, result, q_out );
  input [27:0] divided;
  input [19:0] divisor;
  input [7:0] q_in;
  output [19:0] divisor_out;
  output [27:0] result;
  output [7:0] q_out;
  input clock, reset_n, start;
  output start_out;
  wire   N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N75,
         N76, N77, N78, N79, N80, N81, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313;
  wire   [20:0] stage_result;

  DFFR_X1 start_out_reg ( .D(n229), .CK(clock), .RN(n234), .Q(start_out) );
  DFFR_X1 \q_out_reg[7]  ( .D(N81), .CK(clock), .RN(n234), .Q(q_out[7]) );
  DFFR_X1 \q_out_reg[6]  ( .D(N80), .CK(clock), .RN(n234), .Q(q_out[6]) );
  DFFR_X1 \q_out_reg[5]  ( .D(N79), .CK(clock), .RN(n234), .Q(q_out[5]) );
  DFFR_X1 \q_out_reg[4]  ( .D(N78), .CK(clock), .RN(n234), .Q(q_out[4]) );
  DFFR_X1 \q_out_reg[3]  ( .D(N77), .CK(clock), .RN(n234), .Q(q_out[3]) );
  DFFR_X1 \q_out_reg[2]  ( .D(N76), .CK(clock), .RN(n234), .Q(q_out[2]) );
  DFFR_X1 \q_out_reg[1]  ( .D(N75), .CK(clock), .RN(n234), .Q(q_out[1]) );
  DFFR_X1 \q_out_reg[0]  ( .D(n293), .CK(clock), .RN(n233), .Q(q_out[0]) );
  DFFR_X1 \result_reg[27]  ( .D(n313), .CK(clock), .RN(n233), .Q(result[27])
         );
  DFFR_X1 \result_reg[26]  ( .D(n312), .CK(clock), .RN(n233), .Q(result[26])
         );
  DFFR_X1 \result_reg[25]  ( .D(n311), .CK(clock), .RN(n233), .Q(result[25])
         );
  DFFR_X1 \result_reg[24]  ( .D(n310), .CK(clock), .RN(n233), .Q(result[24])
         );
  DFFR_X1 \result_reg[23]  ( .D(n309), .CK(clock), .RN(n233), .Q(result[23])
         );
  DFFR_X1 \result_reg[22]  ( .D(n308), .CK(clock), .RN(n233), .Q(result[22])
         );
  DFFR_X1 \result_reg[21]  ( .D(n307), .CK(clock), .RN(n233), .Q(result[21])
         );
  DFFR_X1 \result_reg[20]  ( .D(n306), .CK(clock), .RN(n233), .Q(result[20])
         );
  DFFR_X1 \result_reg[19]  ( .D(n305), .CK(clock), .RN(n233), .Q(result[19])
         );
  DFFR_X1 \result_reg[18]  ( .D(n304), .CK(clock), .RN(n233), .Q(result[18])
         );
  DFFR_X1 \result_reg[17]  ( .D(n303), .CK(clock), .RN(n233), .Q(result[17])
         );
  DFFR_X1 \result_reg[16]  ( .D(n302), .CK(clock), .RN(n232), .Q(result[16])
         );
  DFFR_X1 \result_reg[15]  ( .D(n301), .CK(clock), .RN(n232), .Q(result[15])
         );
  DFFR_X1 \result_reg[14]  ( .D(n300), .CK(clock), .RN(n232), .Q(result[14])
         );
  DFFR_X1 \result_reg[13]  ( .D(n299), .CK(clock), .RN(n232), .Q(result[13])
         );
  DFFR_X1 \result_reg[12]  ( .D(n298), .CK(clock), .RN(n232), .Q(result[12])
         );
  DFFR_X1 \result_reg[11]  ( .D(n297), .CK(clock), .RN(n232), .Q(result[11])
         );
  DFFR_X1 \result_reg[10]  ( .D(n296), .CK(clock), .RN(n232), .Q(result[10])
         );
  DFFR_X1 \result_reg[9]  ( .D(n295), .CK(clock), .RN(n232), .Q(result[9]) );
  DFFR_X1 \result_reg[8]  ( .D(n294), .CK(clock), .RN(n232), .Q(result[8]) );
  DFFR_X1 \result_reg[7]  ( .D(N53), .CK(clock), .RN(n232), .Q(result[7]) );
  DFFR_X1 \result_reg[6]  ( .D(N52), .CK(clock), .RN(n232), .Q(result[6]) );
  DFFR_X1 \result_reg[5]  ( .D(N51), .CK(clock), .RN(n232), .Q(result[5]) );
  DFFR_X1 \result_reg[4]  ( .D(N50), .CK(clock), .RN(n233), .Q(result[4]) );
  DFFR_X1 \result_reg[3]  ( .D(N49), .CK(clock), .RN(n231), .Q(result[3]) );
  DFFR_X1 \result_reg[2]  ( .D(N48), .CK(clock), .RN(n234), .Q(result[2]) );
  DFFR_X1 \result_reg[1]  ( .D(N47), .CK(clock), .RN(n234), .Q(result[1]) );
  DFFR_X1 \divisor_out_reg[19]  ( .D(N46), .CK(clock), .RN(n233), .Q(
        divisor_out[19]) );
  DFFR_X1 \divisor_out_reg[18]  ( .D(N45), .CK(clock), .RN(n232), .Q(
        divisor_out[18]) );
  DFFR_X1 \divisor_out_reg[17]  ( .D(N44), .CK(clock), .RN(n231), .Q(
        divisor_out[17]) );
  DFFR_X1 \divisor_out_reg[16]  ( .D(N43), .CK(clock), .RN(n234), .Q(
        divisor_out[16]) );
  DFFR_X1 \divisor_out_reg[15]  ( .D(N42), .CK(clock), .RN(n231), .Q(
        divisor_out[15]) );
  DFFR_X1 \divisor_out_reg[14]  ( .D(N41), .CK(clock), .RN(n234), .Q(
        divisor_out[14]) );
  DFFR_X1 \divisor_out_reg[13]  ( .D(N40), .CK(clock), .RN(n232), .Q(
        divisor_out[13]) );
  DFFR_X1 \divisor_out_reg[12]  ( .D(N39), .CK(clock), .RN(n234), .Q(
        divisor_out[12]) );
  DFFR_X1 \divisor_out_reg[11]  ( .D(N38), .CK(clock), .RN(n231), .Q(
        divisor_out[11]) );
  DFFR_X1 \divisor_out_reg[10]  ( .D(N37), .CK(clock), .RN(n231), .Q(
        divisor_out[10]) );
  DFFR_X1 \divisor_out_reg[9]  ( .D(N36), .CK(clock), .RN(n231), .Q(
        divisor_out[9]) );
  DFFR_X1 \divisor_out_reg[8]  ( .D(N35), .CK(clock), .RN(n231), .Q(
        divisor_out[8]) );
  DFFR_X1 \divisor_out_reg[7]  ( .D(N34), .CK(clock), .RN(n231), .Q(
        divisor_out[7]) );
  DFFR_X1 \divisor_out_reg[6]  ( .D(N33), .CK(clock), .RN(n231), .Q(
        divisor_out[6]) );
  DFFR_X1 \divisor_out_reg[5]  ( .D(N32), .CK(clock), .RN(n231), .Q(
        divisor_out[5]) );
  DFFR_X1 \divisor_out_reg[4]  ( .D(N31), .CK(clock), .RN(n231), .Q(
        divisor_out[4]) );
  DFFR_X1 \divisor_out_reg[3]  ( .D(N30), .CK(clock), .RN(n231), .Q(
        divisor_out[3]) );
  DFFR_X1 \divisor_out_reg[2]  ( .D(N29), .CK(clock), .RN(n231), .Q(
        divisor_out[2]) );
  DFFR_X1 \divisor_out_reg[1]  ( .D(N28), .CK(clock), .RN(n231), .Q(
        divisor_out[1]) );
  DFFR_X1 \divisor_out_reg[0]  ( .D(N27), .CK(clock), .RN(n231), .Q(
        divisor_out[0]) );
  AND2_X1 U47 ( .A1(n229), .A2(q_in[6]), .ZN(N81) );
  AND2_X1 U48 ( .A1(q_in[5]), .A2(n229), .ZN(N80) );
  AND2_X1 U49 ( .A1(q_in[4]), .A2(n229), .ZN(N79) );
  AND2_X1 U50 ( .A1(q_in[3]), .A2(n229), .ZN(N78) );
  AND2_X1 U51 ( .A1(q_in[2]), .A2(n229), .ZN(N77) );
  AND2_X1 U52 ( .A1(q_in[1]), .A2(n229), .ZN(N76) );
  AND2_X1 U53 ( .A1(q_in[0]), .A2(n229), .ZN(N75) );
  AND2_X1 U56 ( .A1(divided[5]), .A2(n229), .ZN(N52) );
  AND2_X1 U57 ( .A1(divided[4]), .A2(n229), .ZN(N51) );
  AND2_X1 U58 ( .A1(divided[3]), .A2(n229), .ZN(N50) );
  AND2_X1 U59 ( .A1(divided[2]), .A2(n229), .ZN(N49) );
  AND2_X1 U60 ( .A1(divided[1]), .A2(n229), .ZN(N48) );
  AND2_X1 U61 ( .A1(divided[0]), .A2(n229), .ZN(N47) );
  AND2_X1 U62 ( .A1(divisor[19]), .A2(n229), .ZN(N46) );
  AND2_X1 U63 ( .A1(divisor[18]), .A2(n229), .ZN(N45) );
  AND2_X1 U64 ( .A1(divisor[17]), .A2(n229), .ZN(N44) );
  AND2_X1 U65 ( .A1(divisor[16]), .A2(n229), .ZN(N43) );
  AND2_X1 U66 ( .A1(divisor[15]), .A2(n229), .ZN(N42) );
  AND2_X1 U67 ( .A1(divisor[14]), .A2(n229), .ZN(N41) );
  AND2_X1 U68 ( .A1(divisor[13]), .A2(n229), .ZN(N40) );
  divider_pipe_stage_3_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(result[0]) );
  INV_X4 U6 ( .A(n235), .ZN(n232) );
  INV_X4 U7 ( .A(n235), .ZN(n233) );
  INV_X4 U8 ( .A(n235), .ZN(n231) );
  INV_X4 U9 ( .A(n235), .ZN(n234) );
  INV_X4 U10 ( .A(reset_n), .ZN(n235) );
  NAND2_X2 U11 ( .A1(n229), .A2(n236), .ZN(n277) );
  NAND2_X2 U12 ( .A1(n229), .A2(n236), .ZN(n225) );
  NAND2_X2 U13 ( .A1(n229), .A2(n236), .ZN(n226) );
  INV_X4 U14 ( .A(n230), .ZN(n229) );
  INV_X4 U15 ( .A(start), .ZN(n230) );
  NAND2_X2 U16 ( .A1(n229), .A2(n237), .ZN(n227) );
  NAND2_X2 U17 ( .A1(n229), .A2(n237), .ZN(n228) );
  XNOR2_X2 U18 ( .A(divided[27]), .B(stage_result[20]), .ZN(n237) );
  INV_X4 U19 ( .A(n237), .ZN(n236) );
  INV_X4 U20 ( .A(n277), .ZN(n293) );
  AND2_X1 U21 ( .A1(divided[6]), .A2(n229), .ZN(N53) );
  NAND2_X2 U22 ( .A1(n229), .A2(n237), .ZN(n279) );
  INV_X4 U23 ( .A(divided[7]), .ZN(n239) );
  INV_X4 U24 ( .A(stage_result[0]), .ZN(n238) );
  OAI22_X2 U25 ( .A1(n227), .A2(n239), .B1(n225), .B2(n238), .ZN(n294) );
  INV_X4 U26 ( .A(divided[8]), .ZN(n241) );
  INV_X4 U27 ( .A(stage_result[1]), .ZN(n240) );
  OAI22_X2 U28 ( .A1(n228), .A2(n241), .B1(n226), .B2(n240), .ZN(n295) );
  INV_X4 U29 ( .A(divided[9]), .ZN(n243) );
  INV_X4 U30 ( .A(stage_result[2]), .ZN(n242) );
  OAI22_X2 U31 ( .A1(n279), .A2(n243), .B1(n225), .B2(n242), .ZN(n296) );
  INV_X4 U32 ( .A(divided[10]), .ZN(n245) );
  INV_X4 U33 ( .A(stage_result[3]), .ZN(n244) );
  OAI22_X2 U34 ( .A1(n227), .A2(n245), .B1(n226), .B2(n244), .ZN(n297) );
  INV_X4 U35 ( .A(divided[11]), .ZN(n247) );
  INV_X4 U36 ( .A(stage_result[4]), .ZN(n246) );
  OAI22_X2 U37 ( .A1(n228), .A2(n247), .B1(n277), .B2(n246), .ZN(n298) );
  INV_X4 U38 ( .A(divided[12]), .ZN(n249) );
  INV_X4 U39 ( .A(stage_result[5]), .ZN(n248) );
  OAI22_X2 U40 ( .A1(n279), .A2(n249), .B1(n225), .B2(n248), .ZN(n299) );
  INV_X4 U41 ( .A(divided[13]), .ZN(n251) );
  INV_X4 U42 ( .A(stage_result[6]), .ZN(n250) );
  OAI22_X2 U43 ( .A1(n227), .A2(n251), .B1(n226), .B2(n250), .ZN(n300) );
  INV_X4 U44 ( .A(divided[14]), .ZN(n253) );
  INV_X4 U45 ( .A(stage_result[7]), .ZN(n252) );
  OAI22_X2 U46 ( .A1(n228), .A2(n253), .B1(n277), .B2(n252), .ZN(n301) );
  INV_X4 U54 ( .A(divided[15]), .ZN(n255) );
  INV_X4 U55 ( .A(stage_result[8]), .ZN(n254) );
  OAI22_X2 U69 ( .A1(n279), .A2(n255), .B1(n225), .B2(n254), .ZN(n302) );
  INV_X4 U70 ( .A(divided[16]), .ZN(n257) );
  INV_X4 U71 ( .A(stage_result[9]), .ZN(n256) );
  OAI22_X2 U72 ( .A1(n227), .A2(n257), .B1(n226), .B2(n256), .ZN(n303) );
  INV_X4 U73 ( .A(divided[17]), .ZN(n259) );
  INV_X4 U74 ( .A(stage_result[10]), .ZN(n258) );
  OAI22_X2 U75 ( .A1(n228), .A2(n259), .B1(n277), .B2(n258), .ZN(n304) );
  INV_X4 U76 ( .A(divided[18]), .ZN(n261) );
  INV_X4 U77 ( .A(stage_result[11]), .ZN(n260) );
  OAI22_X2 U78 ( .A1(n279), .A2(n261), .B1(n225), .B2(n260), .ZN(n305) );
  INV_X4 U79 ( .A(divided[19]), .ZN(n263) );
  INV_X4 U80 ( .A(stage_result[12]), .ZN(n262) );
  OAI22_X2 U81 ( .A1(n227), .A2(n263), .B1(n226), .B2(n262), .ZN(n306) );
  INV_X4 U82 ( .A(divided[20]), .ZN(n265) );
  INV_X4 U83 ( .A(stage_result[13]), .ZN(n264) );
  OAI22_X2 U84 ( .A1(n228), .A2(n265), .B1(n277), .B2(n264), .ZN(n307) );
  INV_X4 U85 ( .A(divided[21]), .ZN(n267) );
  INV_X4 U86 ( .A(stage_result[14]), .ZN(n266) );
  OAI22_X2 U87 ( .A1(n279), .A2(n267), .B1(n225), .B2(n266), .ZN(n308) );
  INV_X4 U88 ( .A(divided[22]), .ZN(n269) );
  INV_X4 U89 ( .A(stage_result[15]), .ZN(n268) );
  OAI22_X2 U90 ( .A1(n227), .A2(n269), .B1(n226), .B2(n268), .ZN(n309) );
  INV_X4 U91 ( .A(divided[23]), .ZN(n271) );
  INV_X4 U92 ( .A(stage_result[16]), .ZN(n270) );
  OAI22_X2 U93 ( .A1(n228), .A2(n271), .B1(n277), .B2(n270), .ZN(n310) );
  INV_X4 U94 ( .A(divided[24]), .ZN(n273) );
  INV_X4 U95 ( .A(stage_result[17]), .ZN(n272) );
  OAI22_X2 U96 ( .A1(n279), .A2(n273), .B1(n225), .B2(n272), .ZN(n311) );
  INV_X4 U97 ( .A(divided[25]), .ZN(n275) );
  INV_X4 U98 ( .A(stage_result[18]), .ZN(n274) );
  OAI22_X2 U99 ( .A1(n227), .A2(n275), .B1(n226), .B2(n274), .ZN(n312) );
  INV_X4 U100 ( .A(divided[26]), .ZN(n278) );
  INV_X4 U101 ( .A(stage_result[19]), .ZN(n276) );
  OAI22_X2 U102 ( .A1(n228), .A2(n278), .B1(n277), .B2(n276), .ZN(n313) );
  INV_X4 U103 ( .A(divisor[0]), .ZN(n280) );
  NOR2_X2 U104 ( .A1(n230), .A2(n280), .ZN(N27) );
  INV_X4 U105 ( .A(divisor[1]), .ZN(n281) );
  NOR2_X2 U106 ( .A1(n230), .A2(n281), .ZN(N28) );
  INV_X4 U107 ( .A(divisor[2]), .ZN(n282) );
  NOR2_X2 U108 ( .A1(n230), .A2(n282), .ZN(N29) );
  INV_X4 U109 ( .A(divisor[3]), .ZN(n283) );
  NOR2_X2 U110 ( .A1(n230), .A2(n283), .ZN(N30) );
  INV_X4 U111 ( .A(divisor[4]), .ZN(n284) );
  NOR2_X2 U112 ( .A1(n230), .A2(n284), .ZN(N31) );
  INV_X4 U113 ( .A(divisor[5]), .ZN(n285) );
  NOR2_X2 U114 ( .A1(n230), .A2(n285), .ZN(N32) );
  INV_X4 U115 ( .A(divisor[6]), .ZN(n286) );
  NOR2_X2 U116 ( .A1(n230), .A2(n286), .ZN(N33) );
  INV_X4 U117 ( .A(divisor[7]), .ZN(n287) );
  NOR2_X2 U118 ( .A1(n230), .A2(n287), .ZN(N34) );
  INV_X4 U119 ( .A(divisor[8]), .ZN(n288) );
  NOR2_X2 U120 ( .A1(n230), .A2(n288), .ZN(N35) );
  INV_X4 U121 ( .A(divisor[9]), .ZN(n289) );
  NOR2_X2 U122 ( .A1(n230), .A2(n289), .ZN(N36) );
  INV_X4 U123 ( .A(divisor[10]), .ZN(n290) );
  NOR2_X2 U124 ( .A1(n230), .A2(n290), .ZN(N37) );
  INV_X4 U125 ( .A(divisor[11]), .ZN(n291) );
  NOR2_X2 U126 ( .A1(n230), .A2(n291), .ZN(N38) );
  INV_X4 U127 ( .A(divisor[12]), .ZN(n292) );
  NOR2_X2 U128 ( .A1(n230), .A2(n292), .ZN(N39) );
endmodule


module divider_pipe_stage_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n110, n112, n114,
         n115, n116, n117, n118, n120, n121, n122;

  FA_X1 U2 ( .A(A[19]), .B(B[19]), .CI(n18), .CO(CO), .S(SUM[19]) );
  FA_X1 U3 ( .A(A[18]), .B(B[18]), .CI(n19), .CO(n18), .S(SUM[18]) );
  FA_X1 U4 ( .A(A[17]), .B(B[17]), .CI(n20), .CO(n19), .S(SUM[17]) );
  XOR2_X2 U5 ( .A(n1), .B(n23), .Z(SUM[16]) );
  NAND2_X2 U7 ( .A1(n107), .A2(n22), .ZN(n1) );
  NAND2_X2 U10 ( .A1(A[16]), .A2(B[16]), .ZN(n22) );
  XOR2_X2 U11 ( .A(n2), .B(n32), .Z(SUM[15]) );
  NAND2_X2 U15 ( .A1(n40), .A2(n28), .ZN(n26) );
  NAND2_X2 U19 ( .A1(n108), .A2(n31), .ZN(n2) );
  NAND2_X2 U22 ( .A1(A[15]), .A2(B[15]), .ZN(n31) );
  XNOR2_X2 U23 ( .A(n37), .B(n3), .ZN(SUM[14]) );
  NAND2_X2 U27 ( .A1(n33), .A2(n36), .ZN(n3) );
  NAND2_X2 U30 ( .A1(A[14]), .A2(B[14]), .ZN(n36) );
  XOR2_X2 U31 ( .A(n4), .B(n44), .Z(SUM[13]) );
  NAND2_X2 U37 ( .A1(n110), .A2(n43), .ZN(n4) );
  NAND2_X2 U40 ( .A1(A[13]), .A2(B[13]), .ZN(n43) );
  XOR2_X2 U41 ( .A(n5), .B(n49), .Z(SUM[12]) );
  NAND2_X2 U45 ( .A1(n45), .A2(n48), .ZN(n5) );
  NAND2_X2 U48 ( .A1(A[12]), .A2(B[12]), .ZN(n48) );
  XOR2_X2 U49 ( .A(n6), .B(n57), .Z(SUM[11]) );
  NAND2_X2 U52 ( .A1(n65), .A2(n53), .ZN(n51) );
  NAND2_X2 U56 ( .A1(n112), .A2(n56), .ZN(n6) );
  NAND2_X2 U59 ( .A1(A[11]), .A2(B[11]), .ZN(n56) );
  XNOR2_X2 U60 ( .A(n62), .B(n7), .ZN(SUM[10]) );
  NAND2_X2 U64 ( .A1(n58), .A2(n61), .ZN(n7) );
  NAND2_X2 U67 ( .A1(A[10]), .A2(B[10]), .ZN(n61) );
  XNOR2_X2 U68 ( .A(n69), .B(n8), .ZN(SUM[9]) );
  NAND2_X2 U74 ( .A1(n114), .A2(n68), .ZN(n8) );
  NAND2_X2 U77 ( .A1(A[9]), .A2(B[9]), .ZN(n68) );
  XOR2_X2 U78 ( .A(n9), .B(n72), .Z(SUM[8]) );
  NAND2_X2 U80 ( .A1(n115), .A2(n71), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[8]), .A2(B[8]), .ZN(n71) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[7]) );
  NAND2_X2 U87 ( .A1(n84), .A2(n76), .ZN(n74) );
  NAND2_X2 U91 ( .A1(n116), .A2(n79), .ZN(n10) );
  NAND2_X2 U94 ( .A1(A[7]), .A2(B[7]), .ZN(n79) );
  XOR2_X2 U95 ( .A(n11), .B(n83), .Z(SUM[6]) );
  NAND2_X2 U97 ( .A1(n117), .A2(n82), .ZN(n11) );
  NAND2_X2 U100 ( .A1(A[6]), .A2(B[6]), .ZN(n82) );
  XOR2_X2 U101 ( .A(n12), .B(n88), .Z(SUM[5]) );
  NAND2_X2 U105 ( .A1(n118), .A2(n87), .ZN(n12) );
  NAND2_X2 U108 ( .A1(A[5]), .A2(B[5]), .ZN(n87) );
  XNOR2_X2 U109 ( .A(n93), .B(n13), .ZN(SUM[4]) );
  NAND2_X2 U113 ( .A1(n89), .A2(n92), .ZN(n13) );
  NAND2_X2 U116 ( .A1(A[4]), .A2(B[4]), .ZN(n92) );
  XNOR2_X2 U117 ( .A(n99), .B(n14), .ZN(SUM[3]) );
  NAND2_X2 U122 ( .A1(n120), .A2(n98), .ZN(n14) );
  NAND2_X2 U125 ( .A1(A[3]), .A2(B[3]), .ZN(n98) );
  XOR2_X2 U126 ( .A(n15), .B(n102), .Z(SUM[2]) );
  NAND2_X2 U128 ( .A1(n121), .A2(n101), .ZN(n15) );
  NAND2_X2 U131 ( .A1(A[2]), .A2(B[2]), .ZN(n101) );
  XOR2_X2 U132 ( .A(n106), .B(n16), .Z(SUM[1]) );
  NAND2_X2 U135 ( .A1(n122), .A2(n105), .ZN(n16) );
  NAND2_X2 U138 ( .A1(A[1]), .A2(B[1]), .ZN(n105) );
  XNOR2_X2 U139 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U144 ( .B1(n73), .B2(n24), .A(n25), .ZN(n23) );
  NOR2_X2 U145 ( .A1(n51), .A2(n26), .ZN(n24) );
  OAI21_X2 U146 ( .B1(n52), .B2(n26), .A(n27), .ZN(n25) );
  OAI21_X2 U147 ( .B1(n49), .B2(n38), .A(n39), .ZN(n37) );
  OAI21_X2 U148 ( .B1(n72), .B2(n51), .A(n52), .ZN(n50) );
  AOI21_X2 U149 ( .B1(n93), .B2(n84), .A(n85), .ZN(n83) );
  OAI21_X2 U150 ( .B1(n72), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X2 U151 ( .B1(n53), .B2(n66), .A(n54), .ZN(n52) );
  OAI21_X2 U152 ( .B1(n55), .B2(n61), .A(n56), .ZN(n54) );
  AOI21_X2 U153 ( .B1(n95), .B2(n103), .A(n96), .ZN(n94) );
  NOR2_X2 U154 ( .A1(n100), .A2(n97), .ZN(n95) );
  OAI21_X2 U155 ( .B1(n97), .B2(n101), .A(n98), .ZN(n96) );
  OAI21_X2 U156 ( .B1(n86), .B2(n92), .A(n87), .ZN(n85) );
  OAI21_X2 U157 ( .B1(n94), .B2(n74), .A(n75), .ZN(n73) );
  AOI21_X2 U158 ( .B1(n76), .B2(n85), .A(n77), .ZN(n75) );
  NOR2_X2 U159 ( .A1(n81), .A2(n78), .ZN(n76) );
  AOI21_X2 U160 ( .B1(n28), .B2(n41), .A(n29), .ZN(n27) );
  OAI21_X2 U161 ( .B1(n30), .B2(n36), .A(n31), .ZN(n29) );
  OAI21_X2 U162 ( .B1(n42), .B2(n48), .A(n43), .ZN(n41) );
  OAI21_X2 U163 ( .B1(n104), .B2(n106), .A(n105), .ZN(n103) );
  OAI21_X2 U164 ( .B1(n67), .B2(n71), .A(n68), .ZN(n66) );
  OAI21_X2 U165 ( .B1(n78), .B2(n82), .A(n79), .ZN(n77) );
  NOR2_X2 U166 ( .A1(n60), .A2(n55), .ZN(n53) );
  NOR2_X2 U167 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U168 ( .A1(n91), .A2(n86), .ZN(n84) );
  NOR2_X2 U169 ( .A1(n70), .A2(n67), .ZN(n65) );
  NOR2_X2 U170 ( .A1(n47), .A2(n42), .ZN(n40) );
  AOI21_X2 U171 ( .B1(n37), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U172 ( .B1(n93), .B2(n89), .A(n90), .ZN(n88) );
  AOI21_X2 U173 ( .B1(n62), .B2(n58), .A(n59), .ZN(n57) );
  AOI21_X2 U174 ( .B1(n50), .B2(n45), .A(n46), .ZN(n44) );
  OAI21_X2 U175 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X2 U176 ( .B1(n83), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U177 ( .B1(n72), .B2(n70), .A(n71), .ZN(n69) );
  OAI21_X2 U178 ( .B1(n23), .B2(n21), .A(n22), .ZN(n20) );
  NOR2_X2 U179 ( .A1(A[3]), .A2(B[3]), .ZN(n97) );
  NOR2_X2 U180 ( .A1(A[7]), .A2(B[7]), .ZN(n78) );
  NOR2_X2 U181 ( .A1(A[5]), .A2(B[5]), .ZN(n86) );
  NOR2_X2 U182 ( .A1(A[11]), .A2(B[11]), .ZN(n55) );
  NOR2_X2 U183 ( .A1(A[9]), .A2(B[9]), .ZN(n67) );
  NOR2_X2 U184 ( .A1(A[15]), .A2(B[15]), .ZN(n30) );
  NOR2_X2 U185 ( .A1(A[13]), .A2(B[13]), .ZN(n42) );
  NOR2_X2 U186 ( .A1(A[2]), .A2(B[2]), .ZN(n100) );
  NOR2_X2 U187 ( .A1(A[6]), .A2(B[6]), .ZN(n81) );
  NOR2_X2 U188 ( .A1(A[8]), .A2(B[8]), .ZN(n70) );
  NOR2_X2 U189 ( .A1(A[1]), .A2(B[1]), .ZN(n104) );
  NOR2_X2 U190 ( .A1(A[0]), .A2(B[0]), .ZN(n106) );
  NOR2_X2 U191 ( .A1(A[4]), .A2(B[4]), .ZN(n91) );
  NOR2_X2 U192 ( .A1(A[10]), .A2(B[10]), .ZN(n60) );
  NOR2_X2 U193 ( .A1(A[12]), .A2(B[12]), .ZN(n47) );
  NOR2_X2 U194 ( .A1(A[14]), .A2(B[14]), .ZN(n35) );
  NOR2_X2 U195 ( .A1(A[16]), .A2(B[16]), .ZN(n21) );
  INV_X4 U196 ( .A(n94), .ZN(n93) );
  INV_X4 U197 ( .A(n92), .ZN(n90) );
  INV_X4 U198 ( .A(n73), .ZN(n72) );
  INV_X4 U199 ( .A(n66), .ZN(n64) );
  INV_X4 U200 ( .A(n65), .ZN(n63) );
  INV_X4 U201 ( .A(n61), .ZN(n59) );
  INV_X4 U202 ( .A(n50), .ZN(n49) );
  INV_X4 U203 ( .A(n48), .ZN(n46) );
  INV_X4 U204 ( .A(n41), .ZN(n39) );
  INV_X4 U205 ( .A(n40), .ZN(n38) );
  INV_X4 U206 ( .A(n36), .ZN(n34) );
  INV_X4 U207 ( .A(n104), .ZN(n122) );
  INV_X4 U208 ( .A(n100), .ZN(n121) );
  INV_X4 U209 ( .A(n97), .ZN(n120) );
  INV_X4 U210 ( .A(n91), .ZN(n89) );
  INV_X4 U211 ( .A(n86), .ZN(n118) );
  INV_X4 U212 ( .A(n81), .ZN(n117) );
  INV_X4 U213 ( .A(n78), .ZN(n116) );
  INV_X4 U214 ( .A(n70), .ZN(n115) );
  INV_X4 U215 ( .A(n67), .ZN(n114) );
  INV_X4 U216 ( .A(n60), .ZN(n58) );
  INV_X4 U217 ( .A(n55), .ZN(n112) );
  INV_X4 U218 ( .A(n47), .ZN(n45) );
  INV_X4 U219 ( .A(n42), .ZN(n110) );
  INV_X4 U220 ( .A(n35), .ZN(n33) );
  INV_X4 U221 ( .A(n30), .ZN(n108) );
  INV_X4 U222 ( .A(n21), .ZN(n107) );
  INV_X4 U223 ( .A(n103), .ZN(n102) );
endmodule


module divider_pipe_stage_2 ( clock, reset_n, start, divided, divisor, q_in, 
        start_out, divisor_out, result, q_out );
  input [27:0] divided;
  input [19:0] divisor;
  input [7:0] q_in;
  output [19:0] divisor_out;
  output [27:0] result;
  output [7:0] q_out;
  input clock, reset_n, start;
  output start_out;
  wire   N27, N28, N29, N31, N32, N33, N34, N35, N36, N37, N38, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N75, N76, N77,
         N78, N79, N80, N81, n227, n229, n231, n234, n236, n238, n240, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328;
  wire   [20:0] stage_result;

  DFFR_X1 start_out_reg ( .D(n246), .CK(clock), .RN(n250), .Q(start_out) );
  DFFR_X1 \q_out_reg[7]  ( .D(N81), .CK(clock), .RN(n250), .Q(q_out[7]) );
  DFFR_X1 \q_out_reg[6]  ( .D(N80), .CK(clock), .RN(n252), .Q(q_out[6]) );
  DFFR_X1 \q_out_reg[5]  ( .D(N79), .CK(clock), .RN(n251), .Q(q_out[5]) );
  DFFR_X1 \q_out_reg[4]  ( .D(N78), .CK(clock), .RN(n249), .Q(q_out[4]) );
  DFFR_X1 \q_out_reg[3]  ( .D(N77), .CK(clock), .RN(n250), .Q(q_out[3]) );
  DFFR_X1 \q_out_reg[2]  ( .D(N76), .CK(clock), .RN(n252), .Q(q_out[2]) );
  DFFR_X1 \q_out_reg[1]  ( .D(N75), .CK(clock), .RN(n249), .Q(q_out[1]) );
  DFFR_X1 \q_out_reg[0]  ( .D(n308), .CK(clock), .RN(n252), .Q(q_out[0]) );
  DFFR_X1 \result_reg[27]  ( .D(n328), .CK(clock), .RN(n252), .Q(result[27])
         );
  DFFR_X1 \result_reg[26]  ( .D(n327), .CK(clock), .RN(n252), .Q(result[26])
         );
  DFFR_X1 \result_reg[25]  ( .D(n326), .CK(clock), .RN(n252), .Q(result[25])
         );
  DFFR_X1 \result_reg[24]  ( .D(n325), .CK(clock), .RN(n252), .Q(result[24])
         );
  DFFR_X1 \result_reg[23]  ( .D(n324), .CK(clock), .RN(n252), .Q(result[23])
         );
  DFFR_X1 \result_reg[22]  ( .D(n323), .CK(clock), .RN(n252), .Q(result[22])
         );
  DFFR_X1 \result_reg[21]  ( .D(n322), .CK(clock), .RN(n252), .Q(result[21])
         );
  DFFR_X1 \result_reg[20]  ( .D(n321), .CK(clock), .RN(n252), .Q(result[20])
         );
  DFFR_X1 \result_reg[19]  ( .D(n320), .CK(clock), .RN(n252), .Q(result[19])
         );
  DFFR_X1 \result_reg[18]  ( .D(n319), .CK(clock), .RN(n252), .Q(result[18])
         );
  DFFR_X1 \result_reg[17]  ( .D(n318), .CK(clock), .RN(n252), .Q(result[17])
         );
  DFFR_X1 \result_reg[16]  ( .D(n317), .CK(clock), .RN(n251), .Q(result[16])
         );
  DFFR_X1 \result_reg[15]  ( .D(n316), .CK(clock), .RN(n251), .Q(result[15])
         );
  DFFR_X1 \result_reg[14]  ( .D(n315), .CK(clock), .RN(n251), .Q(result[14])
         );
  DFFR_X1 \result_reg[13]  ( .D(n314), .CK(clock), .RN(n251), .Q(result[13])
         );
  DFFR_X1 \result_reg[12]  ( .D(n313), .CK(clock), .RN(n251), .Q(result[12])
         );
  DFFR_X1 \result_reg[11]  ( .D(n312), .CK(clock), .RN(n251), .Q(result[11])
         );
  DFFR_X1 \result_reg[6]  ( .D(N52), .CK(clock), .RN(n251), .Q(result[6]) );
  DFFR_X1 \result_reg[5]  ( .D(N51), .CK(clock), .RN(n251), .Q(result[5]) );
  DFFR_X1 \result_reg[4]  ( .D(N50), .CK(clock), .RN(n250), .Q(result[4]) );
  DFFR_X1 \result_reg[3]  ( .D(N49), .CK(clock), .RN(n250), .Q(result[3]) );
  DFFR_X1 \result_reg[2]  ( .D(N48), .CK(clock), .RN(n250), .Q(result[2]) );
  DFFR_X1 \result_reg[1]  ( .D(N47), .CK(clock), .RN(n250), .Q(result[1]) );
  DFFR_X1 \divisor_out_reg[19]  ( .D(N46), .CK(clock), .RN(n250), .Q(
        divisor_out[19]) );
  DFFR_X1 \divisor_out_reg[18]  ( .D(N45), .CK(clock), .RN(n250), .Q(
        divisor_out[18]) );
  DFFR_X1 \divisor_out_reg[17]  ( .D(N44), .CK(clock), .RN(n250), .Q(
        divisor_out[17]) );
  DFFR_X1 \divisor_out_reg[16]  ( .D(N43), .CK(clock), .RN(n250), .Q(
        divisor_out[16]) );
  DFFR_X1 \divisor_out_reg[15]  ( .D(N42), .CK(clock), .RN(n250), .Q(
        divisor_out[15]) );
  DFFR_X1 \divisor_out_reg[14]  ( .D(N41), .CK(clock), .RN(n250), .Q(
        divisor_out[14]) );
  DFFR_X1 \divisor_out_reg[13]  ( .D(N40), .CK(clock), .RN(n250), .Q(
        divisor_out[13]) );
  DFFR_X1 \divisor_out_reg[11]  ( .D(N38), .CK(clock), .RN(n249), .Q(
        divisor_out[11]) );
  DFFR_X1 \divisor_out_reg[10]  ( .D(N37), .CK(clock), .RN(n249), .Q(
        divisor_out[10]) );
  DFFR_X1 \divisor_out_reg[9]  ( .D(N36), .CK(clock), .RN(n249), .Q(
        divisor_out[9]) );
  DFFR_X1 \divisor_out_reg[8]  ( .D(N35), .CK(clock), .RN(n249), .Q(
        divisor_out[8]) );
  DFFR_X1 \divisor_out_reg[7]  ( .D(N34), .CK(clock), .RN(n249), .Q(
        divisor_out[7]) );
  DFFR_X1 \divisor_out_reg[6]  ( .D(N33), .CK(clock), .RN(n249), .Q(
        divisor_out[6]) );
  DFFR_X1 \divisor_out_reg[5]  ( .D(N32), .CK(clock), .RN(n249), .Q(
        divisor_out[5]) );
  DFFR_X1 \divisor_out_reg[4]  ( .D(N31), .CK(clock), .RN(n249), .Q(
        divisor_out[4]) );
  AND2_X1 U47 ( .A1(n246), .A2(q_in[6]), .ZN(N81) );
  AND2_X1 U48 ( .A1(q_in[5]), .A2(n246), .ZN(N80) );
  AND2_X1 U49 ( .A1(q_in[4]), .A2(n246), .ZN(N79) );
  AND2_X1 U50 ( .A1(q_in[3]), .A2(n246), .ZN(N78) );
  AND2_X1 U51 ( .A1(q_in[2]), .A2(n246), .ZN(N77) );
  AND2_X1 U52 ( .A1(q_in[1]), .A2(n246), .ZN(N76) );
  AND2_X1 U53 ( .A1(q_in[0]), .A2(n246), .ZN(N75) );
  AND2_X1 U56 ( .A1(divided[5]), .A2(n246), .ZN(N52) );
  AND2_X1 U57 ( .A1(divided[4]), .A2(n246), .ZN(N51) );
  AND2_X1 U58 ( .A1(divided[3]), .A2(n246), .ZN(N50) );
  AND2_X1 U59 ( .A1(divided[2]), .A2(n246), .ZN(N49) );
  AND2_X1 U60 ( .A1(divided[1]), .A2(n246), .ZN(N48) );
  AND2_X1 U61 ( .A1(divided[0]), .A2(n246), .ZN(N47) );
  AND2_X1 U62 ( .A1(divisor[19]), .A2(n246), .ZN(N46) );
  AND2_X1 U63 ( .A1(divisor[18]), .A2(n246), .ZN(N45) );
  AND2_X1 U64 ( .A1(divisor[17]), .A2(n246), .ZN(N44) );
  AND2_X1 U65 ( .A1(divisor[16]), .A2(n246), .ZN(N43) );
  AND2_X1 U66 ( .A1(divisor[15]), .A2(n246), .ZN(N42) );
  AND2_X1 U67 ( .A1(divisor[14]), .A2(n246), .ZN(N41) );
  AND2_X1 U68 ( .A1(divisor[13]), .A2(n246), .ZN(N40) );
  divider_pipe_stage_2_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  DFFR_X2 \divisor_out_reg[1]  ( .D(N28), .CK(clock), .RN(n249), .QN(n240) );
  DFFR_X2 \divisor_out_reg[0]  ( .D(N27), .CK(clock), .RN(n249), .QN(n238) );
  DFFR_X2 \result_reg[7]  ( .D(N53), .CK(clock), .RN(n251), .QN(n236) );
  DFFR_X2 \result_reg[8]  ( .D(n309), .CK(clock), .RN(n251), .QN(n234) );
  DFFR_X2 \divisor_out_reg[2]  ( .D(N29), .CK(clock), .RN(n249), .QN(n231) );
  DFFR_X2 \result_reg[9]  ( .D(n310), .CK(clock), .RN(n251), .QN(n229) );
  DFFR_X2 \result_reg[10]  ( .D(n311), .CK(clock), .RN(n251), .QN(n227) );
  SDFFR_X1 \divisor_out_reg[3]  ( .D(1'b0), .SI(divisor[3]), .SE(start), .CK(
        clock), .RN(reset_n), .Q(divisor_out[3]) );
  SDFFR_X1 \divisor_out_reg[12]  ( .D(1'b0), .SI(divisor[12]), .SE(start), 
        .CK(clock), .RN(reset_n), .Q(divisor_out[12]) );
  INV_X4 U4 ( .A(1'b1), .ZN(result[0]) );
  INV_X4 U8 ( .A(n248), .ZN(n251) );
  INV_X4 U9 ( .A(n248), .ZN(n249) );
  INV_X4 U10 ( .A(n248), .ZN(n252) );
  INV_X4 U11 ( .A(n248), .ZN(n250) );
  INV_X4 U12 ( .A(reset_n), .ZN(n248) );
  NAND2_X2 U13 ( .A1(n246), .A2(n253), .ZN(n294) );
  NAND2_X2 U14 ( .A1(n246), .A2(n253), .ZN(n242) );
  NAND2_X2 U15 ( .A1(n246), .A2(n253), .ZN(n243) );
  INV_X4 U16 ( .A(n247), .ZN(n246) );
  INV_X4 U17 ( .A(start), .ZN(n247) );
  INV_X2 U18 ( .A(n227), .ZN(result[10]) );
  INV_X2 U19 ( .A(n229), .ZN(result[9]) );
  INV_X2 U20 ( .A(n231), .ZN(divisor_out[2]) );
  INV_X2 U21 ( .A(n234), .ZN(result[8]) );
  INV_X2 U22 ( .A(n236), .ZN(result[7]) );
  INV_X2 U23 ( .A(n238), .ZN(divisor_out[0]) );
  INV_X2 U24 ( .A(n240), .ZN(divisor_out[1]) );
  NAND2_X2 U25 ( .A1(n246), .A2(n254), .ZN(n244) );
  NAND2_X2 U26 ( .A1(n246), .A2(n254), .ZN(n245) );
  XNOR2_X2 U27 ( .A(divided[27]), .B(stage_result[20]), .ZN(n254) );
  INV_X4 U28 ( .A(n254), .ZN(n253) );
  INV_X4 U29 ( .A(n294), .ZN(n308) );
  AND2_X1 U30 ( .A1(divided[6]), .A2(n246), .ZN(N53) );
  NAND2_X2 U31 ( .A1(n246), .A2(n254), .ZN(n296) );
  INV_X4 U32 ( .A(divided[7]), .ZN(n256) );
  INV_X4 U33 ( .A(stage_result[0]), .ZN(n255) );
  OAI22_X2 U34 ( .A1(n244), .A2(n256), .B1(n242), .B2(n255), .ZN(n309) );
  INV_X4 U35 ( .A(divided[8]), .ZN(n258) );
  INV_X4 U36 ( .A(stage_result[1]), .ZN(n257) );
  OAI22_X2 U37 ( .A1(n245), .A2(n258), .B1(n243), .B2(n257), .ZN(n310) );
  INV_X4 U38 ( .A(divided[9]), .ZN(n260) );
  INV_X4 U39 ( .A(stage_result[2]), .ZN(n259) );
  OAI22_X2 U40 ( .A1(n296), .A2(n260), .B1(n242), .B2(n259), .ZN(n311) );
  INV_X4 U41 ( .A(divided[10]), .ZN(n262) );
  INV_X4 U42 ( .A(stage_result[3]), .ZN(n261) );
  OAI22_X2 U43 ( .A1(n244), .A2(n262), .B1(n243), .B2(n261), .ZN(n312) );
  INV_X4 U44 ( .A(divided[11]), .ZN(n264) );
  INV_X4 U45 ( .A(stage_result[4]), .ZN(n263) );
  OAI22_X2 U46 ( .A1(n245), .A2(n264), .B1(n294), .B2(n263), .ZN(n313) );
  INV_X4 U54 ( .A(divided[12]), .ZN(n266) );
  INV_X4 U55 ( .A(stage_result[5]), .ZN(n265) );
  OAI22_X2 U69 ( .A1(n296), .A2(n266), .B1(n242), .B2(n265), .ZN(n314) );
  INV_X4 U70 ( .A(divided[13]), .ZN(n268) );
  INV_X4 U71 ( .A(stage_result[6]), .ZN(n267) );
  OAI22_X2 U72 ( .A1(n244), .A2(n268), .B1(n243), .B2(n267), .ZN(n315) );
  INV_X4 U73 ( .A(divided[14]), .ZN(n270) );
  INV_X4 U74 ( .A(stage_result[7]), .ZN(n269) );
  OAI22_X2 U75 ( .A1(n245), .A2(n270), .B1(n294), .B2(n269), .ZN(n316) );
  INV_X4 U76 ( .A(divided[15]), .ZN(n272) );
  INV_X4 U77 ( .A(stage_result[8]), .ZN(n271) );
  OAI22_X2 U78 ( .A1(n296), .A2(n272), .B1(n242), .B2(n271), .ZN(n317) );
  INV_X4 U79 ( .A(divided[16]), .ZN(n274) );
  INV_X4 U80 ( .A(stage_result[9]), .ZN(n273) );
  OAI22_X2 U81 ( .A1(n244), .A2(n274), .B1(n243), .B2(n273), .ZN(n318) );
  INV_X4 U82 ( .A(divided[17]), .ZN(n276) );
  INV_X4 U83 ( .A(stage_result[10]), .ZN(n275) );
  OAI22_X2 U84 ( .A1(n245), .A2(n276), .B1(n294), .B2(n275), .ZN(n319) );
  INV_X4 U85 ( .A(divided[18]), .ZN(n278) );
  INV_X4 U86 ( .A(stage_result[11]), .ZN(n277) );
  OAI22_X2 U87 ( .A1(n296), .A2(n278), .B1(n242), .B2(n277), .ZN(n320) );
  INV_X4 U88 ( .A(divided[19]), .ZN(n280) );
  INV_X4 U89 ( .A(stage_result[12]), .ZN(n279) );
  OAI22_X2 U90 ( .A1(n244), .A2(n280), .B1(n243), .B2(n279), .ZN(n321) );
  INV_X4 U91 ( .A(divided[20]), .ZN(n282) );
  INV_X4 U92 ( .A(stage_result[13]), .ZN(n281) );
  OAI22_X2 U93 ( .A1(n245), .A2(n282), .B1(n294), .B2(n281), .ZN(n322) );
  INV_X4 U94 ( .A(divided[21]), .ZN(n284) );
  INV_X4 U95 ( .A(stage_result[14]), .ZN(n283) );
  OAI22_X2 U96 ( .A1(n296), .A2(n284), .B1(n242), .B2(n283), .ZN(n323) );
  INV_X4 U97 ( .A(divided[22]), .ZN(n286) );
  INV_X4 U98 ( .A(stage_result[15]), .ZN(n285) );
  OAI22_X2 U99 ( .A1(n244), .A2(n286), .B1(n243), .B2(n285), .ZN(n324) );
  INV_X4 U100 ( .A(divided[23]), .ZN(n288) );
  INV_X4 U101 ( .A(stage_result[16]), .ZN(n287) );
  OAI22_X2 U102 ( .A1(n245), .A2(n288), .B1(n294), .B2(n287), .ZN(n325) );
  INV_X4 U103 ( .A(divided[24]), .ZN(n290) );
  INV_X4 U104 ( .A(stage_result[17]), .ZN(n289) );
  OAI22_X2 U105 ( .A1(n296), .A2(n290), .B1(n242), .B2(n289), .ZN(n326) );
  INV_X4 U106 ( .A(divided[25]), .ZN(n292) );
  INV_X4 U107 ( .A(stage_result[18]), .ZN(n291) );
  OAI22_X2 U108 ( .A1(n244), .A2(n292), .B1(n243), .B2(n291), .ZN(n327) );
  INV_X4 U109 ( .A(divided[26]), .ZN(n295) );
  INV_X4 U110 ( .A(stage_result[19]), .ZN(n293) );
  OAI22_X2 U111 ( .A1(n245), .A2(n295), .B1(n294), .B2(n293), .ZN(n328) );
  INV_X4 U112 ( .A(divisor[0]), .ZN(n297) );
  NOR2_X2 U113 ( .A1(n247), .A2(n297), .ZN(N27) );
  INV_X4 U114 ( .A(divisor[1]), .ZN(n298) );
  NOR2_X2 U115 ( .A1(n247), .A2(n298), .ZN(N28) );
  INV_X4 U116 ( .A(divisor[2]), .ZN(n299) );
  NOR2_X2 U117 ( .A1(n247), .A2(n299), .ZN(N29) );
  INV_X4 U118 ( .A(divisor[4]), .ZN(n300) );
  NOR2_X2 U119 ( .A1(n247), .A2(n300), .ZN(N31) );
  INV_X4 U120 ( .A(divisor[5]), .ZN(n301) );
  NOR2_X2 U121 ( .A1(n247), .A2(n301), .ZN(N32) );
  INV_X4 U122 ( .A(divisor[6]), .ZN(n302) );
  NOR2_X2 U123 ( .A1(n247), .A2(n302), .ZN(N33) );
  INV_X4 U124 ( .A(divisor[7]), .ZN(n303) );
  NOR2_X2 U125 ( .A1(n247), .A2(n303), .ZN(N34) );
  INV_X4 U126 ( .A(divisor[8]), .ZN(n304) );
  NOR2_X2 U127 ( .A1(n247), .A2(n304), .ZN(N35) );
  INV_X4 U128 ( .A(divisor[9]), .ZN(n305) );
  NOR2_X2 U129 ( .A1(n247), .A2(n305), .ZN(N36) );
  INV_X4 U130 ( .A(divisor[10]), .ZN(n306) );
  NOR2_X2 U131 ( .A1(n247), .A2(n306), .ZN(N37) );
  INV_X4 U132 ( .A(divisor[11]), .ZN(n307) );
  NOR2_X2 U133 ( .A1(n247), .A2(n307), .ZN(N38) );
endmodule


module divider_pipe_stage_0 ( clock, reset_n, start, divided, divisor, q_in, 
        start_out, divisor_out, result, q_out );
  input [27:0] divided;
  input [19:0] divisor;
  input [7:0] q_in;
  output [19:0] divisor_out;
  output [27:0] result;
  output [7:0] q_out;
  input clock, reset_n, start;
  output start_out;
  wire   \U7/Z_0 , \U7/Z_1 , \U7/Z_2 , \U7/Z_3 , \U7/Z_4 , \U7/Z_5 , \U7/Z_6 ,
         \U7/Z_7 , \U7/Z_8 , \U7/Z_9 , \U7/Z_10 , \U7/Z_11 , \U7/Z_12 ,
         \U7/Z_13 , \U7/Z_14 , \U7/Z_15 , \U7/Z_16 , \U7/Z_17 , \U7/Z_18 ,
         \U7/Z_19 , \U7/DATA1_0 , \U7/DATA1_1 , \U7/DATA1_2 , \U7/DATA1_3 ,
         \U7/DATA1_4 , \U7/DATA1_5 , \U7/DATA1_6 , \U7/DATA1_7 , \U7/DATA1_8 ,
         \U7/DATA1_9 , \U7/DATA1_10 , \U7/DATA1_11 , \U7/DATA1_12 ,
         \U7/DATA1_13 , \U7/DATA1_14 , \U7/DATA1_15 , \U7/DATA1_16 ,
         \U7/DATA1_17 , \U7/DATA1_18 , \U7/DATA1_19 , \U6/Z_0 , \U6/Z_1 ,
         \U6/Z_2 , \U6/Z_3 , \U6/Z_4 , \U6/Z_5 , \U6/Z_6 , \U6/DATA1_0 ,
         \U6/DATA1_1 , \U6/DATA1_2 , \U6/DATA1_3 , \U6/DATA1_4 , \U6/DATA1_5 ,
         \U6/DATA1_6 , \U5/Z_1 , \U5/Z_2 , \U5/Z_3 , \U5/Z_4 , \U5/Z_5 ,
         \U5/Z_6 , \U5/Z_7 , \U5/DATA1_1 , \U5/DATA1_2 , \U5/DATA1_3 ,
         \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 , \U5/DATA1_7 , \U4/DATA2_0 ,
         \U4/DATA2_1 , \U4/DATA2_2 , \U4/DATA2_3 , \U4/DATA2_4 , \U4/DATA2_5 ,
         \U4/DATA2_6 , \U4/DATA2_7 , \U4/DATA2_8 , \U4/DATA2_9 , \U4/DATA2_10 ,
         \U4/DATA2_11 , \U4/DATA2_12 , \U4/DATA2_13 , \U4/DATA2_14 ,
         \U4/DATA2_15 , \U4/DATA2_16 , \U4/DATA2_17 , \U4/DATA2_18 ,
         \U4/DATA2_19 , n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428;
  assign \U7/DATA1_0  = divisor[0];
  assign \U7/DATA1_1  = divisor[1];
  assign \U7/DATA1_2  = divisor[2];
  assign \U7/DATA1_3  = divisor[3];
  assign \U7/DATA1_4  = divisor[4];
  assign \U7/DATA1_5  = divisor[5];
  assign \U7/DATA1_6  = divisor[6];
  assign \U7/DATA1_7  = divisor[7];
  assign \U7/DATA1_8  = divisor[8];
  assign \U7/DATA1_9  = divisor[9];
  assign \U7/DATA1_10  = divisor[10];
  assign \U7/DATA1_11  = divisor[11];
  assign \U7/DATA1_12  = divisor[12];
  assign \U7/DATA1_13  = divisor[13];
  assign \U7/DATA1_14  = divisor[14];
  assign \U7/DATA1_15  = divisor[15];
  assign \U7/DATA1_16  = divisor[16];
  assign \U7/DATA1_17  = divisor[17];
  assign \U7/DATA1_18  = divisor[18];
  assign \U7/DATA1_19  = divisor[19];
  assign \U6/DATA1_0  = divided[0];
  assign \U6/DATA1_1  = divided[1];
  assign \U6/DATA1_2  = divided[2];
  assign \U6/DATA1_3  = divided[3];
  assign \U6/DATA1_4  = divided[4];
  assign \U6/DATA1_5  = divided[5];
  assign \U6/DATA1_6  = divided[6];
  assign \U5/DATA1_1  = q_in[0];
  assign \U5/DATA1_2  = q_in[1];
  assign \U5/DATA1_3  = q_in[2];
  assign \U5/DATA1_4  = q_in[3];
  assign \U5/DATA1_5  = q_in[4];
  assign \U5/DATA1_6  = q_in[5];
  assign \U5/DATA1_7  = q_in[6];
  assign \U4/DATA2_0  = divided[7];
  assign \U4/DATA2_1  = divided[8];
  assign \U4/DATA2_2  = divided[9];
  assign \U4/DATA2_3  = divided[10];
  assign \U4/DATA2_4  = divided[11];
  assign \U4/DATA2_5  = divided[12];
  assign \U4/DATA2_6  = divided[13];
  assign \U4/DATA2_7  = divided[14];
  assign \U4/DATA2_8  = divided[15];
  assign \U4/DATA2_9  = divided[16];
  assign \U4/DATA2_10  = divided[17];
  assign \U4/DATA2_11  = divided[18];
  assign \U4/DATA2_12  = divided[19];
  assign \U4/DATA2_13  = divided[20];
  assign \U4/DATA2_14  = divided[21];
  assign \U4/DATA2_15  = divided[22];
  assign \U4/DATA2_16  = divided[23];
  assign \U4/DATA2_17  = divided[24];
  assign \U4/DATA2_18  = divided[25];
  assign \U4/DATA2_19  = divided[26];

  DFFR_X1 \q_out_reg[7]  ( .D(\U5/Z_7 ), .CK(clock), .RN(n270), .Q(q_out[7])
         );
  DFFR_X1 \q_out_reg[6]  ( .D(\U5/Z_6 ), .CK(clock), .RN(n270), .Q(q_out[6])
         );
  DFFR_X1 \q_out_reg[5]  ( .D(\U5/Z_5 ), .CK(clock), .RN(n270), .Q(q_out[5])
         );
  DFFR_X1 \q_out_reg[4]  ( .D(\U5/Z_4 ), .CK(clock), .RN(n270), .Q(q_out[4])
         );
  DFFR_X1 \q_out_reg[3]  ( .D(\U5/Z_3 ), .CK(clock), .RN(n270), .Q(q_out[3])
         );
  DFFR_X1 \q_out_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .RN(n270), .Q(q_out[2])
         );
  DFFR_X1 \q_out_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .RN(n270), .Q(q_out[1])
         );
  DFFR_X1 \result_reg[7]  ( .D(\U6/Z_6 ), .CK(clock), .RN(n268), .Q(result[7])
         );
  DFFR_X1 \result_reg[6]  ( .D(\U6/Z_5 ), .CK(clock), .RN(n268), .Q(result[6])
         );
  DFFR_X1 \result_reg[5]  ( .D(\U6/Z_4 ), .CK(clock), .RN(n268), .Q(result[5])
         );
  DFFR_X1 \result_reg[4]  ( .D(\U6/Z_3 ), .CK(clock), .RN(n267), .Q(result[4])
         );
  DFFR_X1 \result_reg[3]  ( .D(\U6/Z_2 ), .CK(clock), .RN(reset_n), .Q(
        result[3]) );
  DFFR_X1 \result_reg[2]  ( .D(\U6/Z_1 ), .CK(clock), .RN(n268), .Q(result[2])
         );
  DFFR_X1 \result_reg[1]  ( .D(\U6/Z_0 ), .CK(clock), .RN(n267), .Q(result[1])
         );
  DFFR_X1 \divisor_out_reg[19]  ( .D(\U7/Z_19 ), .CK(clock), .RN(n270), .Q(
        divisor_out[19]) );
  DFFR_X1 \divisor_out_reg[18]  ( .D(\U7/Z_18 ), .CK(clock), .RN(n270), .Q(
        divisor_out[18]) );
  DFFR_X1 \divisor_out_reg[17]  ( .D(\U7/Z_17 ), .CK(clock), .RN(n270), .Q(
        divisor_out[17]) );
  DFFR_X1 \divisor_out_reg[16]  ( .D(\U7/Z_16 ), .CK(clock), .RN(n268), .Q(
        divisor_out[16]) );
  DFFR_X1 \divisor_out_reg[15]  ( .D(\U7/Z_15 ), .CK(clock), .RN(n270), .Q(
        divisor_out[15]) );
  DFFR_X1 \divisor_out_reg[14]  ( .D(\U7/Z_14 ), .CK(clock), .RN(n269), .Q(
        divisor_out[14]) );
  DFFR_X1 \divisor_out_reg[13]  ( .D(\U7/Z_13 ), .CK(clock), .RN(n270), .Q(
        divisor_out[13]) );
  DFFR_X1 \divisor_out_reg[12]  ( .D(\U7/Z_12 ), .CK(clock), .RN(n269), .Q(
        divisor_out[12]) );
  AND2_X1 U55 ( .A1(\U7/DATA1_19 ), .A2(n264), .ZN(\U7/Z_19 ) );
  AND2_X1 U56 ( .A1(\U7/DATA1_18 ), .A2(n264), .ZN(\U7/Z_18 ) );
  AND2_X1 U57 ( .A1(\U7/DATA1_17 ), .A2(n264), .ZN(\U7/Z_17 ) );
  AND2_X1 U58 ( .A1(\U7/DATA1_16 ), .A2(n264), .ZN(\U7/Z_16 ) );
  AND2_X1 U59 ( .A1(\U7/DATA1_15 ), .A2(n264), .ZN(\U7/Z_15 ) );
  AND2_X1 U60 ( .A1(\U7/DATA1_14 ), .A2(n264), .ZN(\U7/Z_14 ) );
  AND2_X1 U61 ( .A1(\U7/DATA1_13 ), .A2(n264), .ZN(\U7/Z_13 ) );
  AND2_X1 U62 ( .A1(\U7/DATA1_12 ), .A2(n264), .ZN(\U7/Z_12 ) );
  AND2_X1 U68 ( .A1(\U6/DATA1_5 ), .A2(n264), .ZN(\U6/Z_5 ) );
  AND2_X1 U69 ( .A1(\U6/DATA1_4 ), .A2(n264), .ZN(\U6/Z_4 ) );
  AND2_X1 U70 ( .A1(\U6/DATA1_3 ), .A2(n264), .ZN(\U6/Z_3 ) );
  AND2_X1 U71 ( .A1(\U6/DATA1_2 ), .A2(n264), .ZN(\U6/Z_2 ) );
  AND2_X1 U72 ( .A1(\U6/DATA1_1 ), .A2(n264), .ZN(\U6/Z_1 ) );
  AND2_X1 U73 ( .A1(\U6/DATA1_0 ), .A2(n264), .ZN(\U6/Z_0 ) );
  AND2_X1 U74 ( .A1(\U5/DATA1_7 ), .A2(n264), .ZN(\U5/Z_7 ) );
  AND2_X1 U75 ( .A1(\U5/DATA1_6 ), .A2(n264), .ZN(\U5/Z_6 ) );
  AND2_X1 U76 ( .A1(\U5/DATA1_5 ), .A2(n264), .ZN(\U5/Z_5 ) );
  AND2_X1 U77 ( .A1(\U5/DATA1_4 ), .A2(n264), .ZN(\U5/Z_4 ) );
  AND2_X1 U78 ( .A1(\U5/DATA1_3 ), .A2(n264), .ZN(\U5/Z_3 ) );
  AND2_X1 U79 ( .A1(\U5/DATA1_2 ), .A2(n264), .ZN(\U5/Z_2 ) );
  AND2_X1 U80 ( .A1(\U5/DATA1_1 ), .A2(n264), .ZN(\U5/Z_1 ) );
  DFFR_X1 \result_reg[25]  ( .D(n423), .CK(clock), .RN(n269), .Q(result[25])
         );
  DFFR_X1 \result_reg[26]  ( .D(n424), .CK(clock), .RN(n269), .Q(result[26])
         );
  DFFR_X1 \result_reg[24]  ( .D(n422), .CK(clock), .RN(n269), .Q(result[24])
         );
  DFFR_X1 \result_reg[27]  ( .D(n425), .CK(clock), .RN(n269), .Q(result[27])
         );
  DFFR_X1 \result_reg[19]  ( .D(n417), .CK(clock), .RN(n269), .Q(result[19])
         );
  DFFR_X1 \result_reg[17]  ( .D(n415), .CK(clock), .RN(n269), .Q(result[17])
         );
  DFFR_X1 \result_reg[23]  ( .D(n421), .CK(clock), .RN(n269), .Q(result[23])
         );
  DFFR_X1 \result_reg[21]  ( .D(n419), .CK(clock), .RN(n269), .Q(result[21])
         );
  DFFR_X1 \result_reg[22]  ( .D(n420), .CK(clock), .RN(n269), .Q(result[22])
         );
  DFFR_X1 \result_reg[16]  ( .D(n414), .CK(clock), .RN(n268), .Q(result[16])
         );
  DFFR_X1 \result_reg[18]  ( .D(n416), .CK(clock), .RN(n269), .Q(result[18])
         );
  DFFR_X1 \result_reg[20]  ( .D(n418), .CK(clock), .RN(n269), .Q(result[20])
         );
  DFFR_X1 \result_reg[13]  ( .D(n411), .CK(clock), .RN(n268), .Q(result[13])
         );
  DFFR_X1 \result_reg[15]  ( .D(n413), .CK(clock), .RN(n268), .Q(result[15])
         );
  DFFR_X1 \result_reg[14]  ( .D(n412), .CK(clock), .RN(n268), .Q(result[14])
         );
  DFFR_X1 \result_reg[12]  ( .D(n410), .CK(clock), .RN(n268), .Q(result[12])
         );
  DFFR_X1 \result_reg[11]  ( .D(n409), .CK(clock), .RN(reset_n), .Q(result[11]) );
  DFFR_X2 \divisor_out_reg[10]  ( .D(\U7/Z_10 ), .CK(clock), .RN(n267), .Q(
        divisor_out[10]) );
  DFFR_X2 \divisor_out_reg[9]  ( .D(\U7/Z_9 ), .CK(clock), .RN(n267), .Q(
        divisor_out[9]) );
  DFFR_X2 \divisor_out_reg[8]  ( .D(\U7/Z_8 ), .CK(clock), .RN(n267), .Q(
        divisor_out[8]) );
  DFFR_X2 \divisor_out_reg[7]  ( .D(\U7/Z_7 ), .CK(clock), .RN(n267), .Q(
        divisor_out[7]) );
  DFFR_X2 \divisor_out_reg[6]  ( .D(\U7/Z_6 ), .CK(clock), .RN(n267), .Q(
        divisor_out[6]) );
  DFFR_X2 \divisor_out_reg[5]  ( .D(\U7/Z_5 ), .CK(clock), .RN(n267), .Q(
        divisor_out[5]) );
  DFFR_X2 \divisor_out_reg[4]  ( .D(\U7/Z_4 ), .CK(clock), .RN(n267), .Q(
        divisor_out[4]) );
  DFFR_X2 \divisor_out_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .RN(n267), .Q(
        divisor_out[2]) );
  DFFR_X2 \divisor_out_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .RN(n267), .Q(
        divisor_out[3]) );
  DFFR_X2 \divisor_out_reg[11]  ( .D(\U7/Z_11 ), .CK(clock), .RN(n267), .Q(
        divisor_out[11]) );
  DFFR_X2 \divisor_out_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .RN(n267), .Q(
        divisor_out[1]) );
  DFFR_X2 \divisor_out_reg[0]  ( .D(\U7/Z_0 ), .CK(clock), .RN(n267), .Q(
        divisor_out[0]) );
  DFFR_X2 start_out_reg ( .D(start), .CK(clock), .RN(n270), .Q(start_out) );
  DFFR_X2 \q_out_reg[0]  ( .D(n408), .CK(clock), .RN(n269), .Q(q_out[0]) );
  DFFR_X2 \result_reg[9]  ( .D(n427), .CK(clock), .RN(n268), .Q(result[9]) );
  DFFR_X2 \result_reg[10]  ( .D(n428), .CK(clock), .RN(n268), .Q(result[10])
         );
  DFFR_X2 \result_reg[8]  ( .D(n426), .CK(clock), .RN(n268), .Q(result[8]) );
  INV_X4 U4 ( .A(1'b1), .ZN(result[0]) );
  NAND2_X2 U6 ( .A1(n324), .A2(n264), .ZN(n263) );
  OAI21_X2 U7 ( .B1(n388), .B2(n308), .A(n307), .ZN(n391) );
  NAND2_X2 U8 ( .A1(n324), .A2(n264), .ZN(n262) );
  INV_X1 U9 ( .A(n231), .ZN(n379) );
  AOI22_X4 U10 ( .A1(n303), .A2(n231), .B1(\U7/DATA1_13 ), .B2(\U4/DATA2_13 ), 
        .ZN(n381) );
  INV_X1 U11 ( .A(n233), .ZN(n385) );
  INV_X4 U12 ( .A(n309), .ZN(n226) );
  NOR2_X2 U13 ( .A1(n323), .A2(n322), .ZN(n324) );
  NAND2_X2 U14 ( .A1(n258), .A2(n264), .ZN(n260) );
  NAND2_X2 U15 ( .A1(n324), .A2(n264), .ZN(n397) );
  INV_X4 U16 ( .A(n259), .ZN(n258) );
  AND2_X4 U17 ( .A1(n394), .A2(n311), .ZN(n225) );
  NAND2_X2 U18 ( .A1(n295), .A2(n294), .ZN(n297) );
  NAND2_X2 U19 ( .A1(n264), .A2(n258), .ZN(n399) );
  OAI22_X2 U20 ( .A1(n377), .A2(n232), .B1(n280), .B2(n281), .ZN(n231) );
  OAI22_X2 U21 ( .A1(n238), .A2(n367), .B1(n368), .B2(n288), .ZN(n237) );
  OAI22_X2 U22 ( .A1(n234), .A2(n383), .B1(n274), .B2(n275), .ZN(n233) );
  NAND2_X1 U23 ( .A1(n391), .A2(n227), .ZN(n317) );
  NOR2_X2 U24 ( .A1(n226), .A2(n230), .ZN(n227) );
  NAND2_X2 U25 ( .A1(n225), .A2(n228), .ZN(n316) );
  NAND2_X2 U26 ( .A1(n309), .A2(n391), .ZN(n228) );
  NAND2_X1 U27 ( .A1(n309), .A2(n391), .ZN(n229) );
  OR2_X1 U28 ( .A1(divided[27]), .A2(n256), .ZN(n230) );
  INV_X4 U29 ( .A(\U7/DATA1_0 ), .ZN(n401) );
  NAND2_X2 U30 ( .A1(n333), .A2(n403), .ZN(n336) );
  XNOR2_X1 U31 ( .A(n383), .B(n244), .ZN(n384) );
  INV_X1 U32 ( .A(n237), .ZN(n370) );
  AND2_X4 U33 ( .A1(n281), .A2(n280), .ZN(n232) );
  AND2_X4 U34 ( .A1(n275), .A2(n274), .ZN(n234) );
  XNOR2_X2 U35 ( .A(n328), .B(n235), .ZN(n330) );
  XOR2_X1 U36 ( .A(\U7/DATA1_1 ), .B(n329), .Z(n235) );
  XNOR2_X1 U37 ( .A(n372), .B(n247), .ZN(n373) );
  XNOR2_X1 U38 ( .A(n381), .B(n248), .ZN(n382) );
  XNOR2_X1 U39 ( .A(n374), .B(n249), .ZN(n375) );
  XNOR2_X1 U40 ( .A(\U7/DATA1_4 ), .B(\U4/DATA2_4 ), .ZN(n250) );
  XNOR2_X1 U41 ( .A(\U7/DATA1_6 ), .B(\U4/DATA2_6 ), .ZN(n251) );
  XNOR2_X1 U42 ( .A(n391), .B(n236), .ZN(n393) );
  XOR2_X2 U43 ( .A(\U7/DATA1_18 ), .B(\U4/DATA2_18 ), .Z(n236) );
  XNOR2_X1 U44 ( .A(\U7/DATA1_7 ), .B(\U4/DATA2_7 ), .ZN(n252) );
  XNOR2_X1 U45 ( .A(\U7/DATA1_5 ), .B(\U4/DATA2_5 ), .ZN(n253) );
  AND2_X4 U46 ( .A1(n368), .A2(n288), .ZN(n238) );
  NOR2_X1 U47 ( .A1(\U4/DATA2_3 ), .A2(\U7/DATA1_3 ), .ZN(n239) );
  NOR2_X4 U48 ( .A1(n291), .A2(n290), .ZN(n240) );
  INV_X1 U49 ( .A(n336), .ZN(n241) );
  OR3_X4 U50 ( .A1(n240), .A2(n239), .A3(n241), .ZN(n342) );
  INV_X4 U51 ( .A(n266), .ZN(n269) );
  INV_X4 U52 ( .A(n266), .ZN(n267) );
  INV_X4 U53 ( .A(n266), .ZN(n268) );
  INV_X4 U54 ( .A(n266), .ZN(n270) );
  INV_X4 U63 ( .A(reset_n), .ZN(n266) );
  XOR2_X2 U64 ( .A(n335), .B(n242), .Z(n334) );
  XNOR2_X2 U65 ( .A(\U7/DATA1_2 ), .B(\U4/DATA2_2 ), .ZN(n242) );
  INV_X4 U66 ( .A(n319), .ZN(n256) );
  INV_X4 U67 ( .A(n265), .ZN(n264) );
  XNOR2_X2 U81 ( .A(n379), .B(n243), .ZN(n380) );
  XNOR2_X2 U82 ( .A(\U7/DATA1_13 ), .B(\U4/DATA2_13 ), .ZN(n243) );
  XNOR2_X2 U83 ( .A(\U7/DATA1_15 ), .B(\U4/DATA2_15 ), .ZN(n244) );
  XNOR2_X2 U84 ( .A(n385), .B(n245), .ZN(n386) );
  XNOR2_X2 U85 ( .A(\U7/DATA1_16 ), .B(\U4/DATA2_16 ), .ZN(n245) );
  XNOR2_X2 U86 ( .A(n370), .B(n246), .ZN(n371) );
  XNOR2_X2 U87 ( .A(\U7/DATA1_9 ), .B(\U4/DATA2_9 ), .ZN(n246) );
  XNOR2_X2 U88 ( .A(\U7/DATA1_10 ), .B(\U4/DATA2_10 ), .ZN(n247) );
  XNOR2_X2 U89 ( .A(\U7/DATA1_14 ), .B(\U4/DATA2_14 ), .ZN(n248) );
  XNOR2_X2 U90 ( .A(\U7/DATA1_11 ), .B(\U4/DATA2_11 ), .ZN(n249) );
  XOR2_X2 U91 ( .A(n346), .B(n250), .Z(n345) );
  XOR2_X2 U92 ( .A(n359), .B(n251), .Z(n358) );
  XOR2_X2 U93 ( .A(n252), .B(n363), .Z(n365) );
  XOR2_X2 U94 ( .A(n253), .B(n349), .Z(n351) );
  INV_X4 U95 ( .A(start), .ZN(n265) );
  INV_X1 U96 ( .A(\U4/DATA2_3 ), .ZN(n254) );
  INV_X1 U97 ( .A(\U4/DATA2_2 ), .ZN(n333) );
  INV_X1 U98 ( .A(\U7/DATA1_2 ), .ZN(n403) );
  INV_X1 U99 ( .A(\U7/DATA1_3 ), .ZN(n255) );
  INV_X1 U100 ( .A(n325), .ZN(n328) );
  NOR2_X1 U101 ( .A1(n265), .A2(n402), .ZN(\U7/Z_1 ) );
  NAND2_X1 U102 ( .A1(n338), .A2(n337), .ZN(n339) );
  INV_X4 U103 ( .A(\U4/DATA2_0 ), .ZN(n326) );
  NOR2_X1 U104 ( .A1(n265), .A2(n401), .ZN(\U7/Z_0 ) );
  INV_X4 U105 ( .A(\U7/DATA1_1 ), .ZN(n402) );
  INV_X2 U106 ( .A(n399), .ZN(n408) );
  NAND2_X1 U107 ( .A1(n332), .A2(n331), .ZN(n335) );
  INV_X2 U108 ( .A(n331), .ZN(n291) );
  NAND2_X1 U109 ( .A1(\U4/DATA2_3 ), .A2(\U7/DATA1_3 ), .ZN(n343) );
  NAND2_X2 U110 ( .A1(n264), .A2(n258), .ZN(n257) );
  NAND2_X2 U111 ( .A1(n264), .A2(n258), .ZN(n261) );
  XOR2_X1 U112 ( .A(\U7/DATA1_3 ), .B(\U4/DATA2_3 ), .Z(n340) );
  NOR2_X2 U113 ( .A1(n323), .A2(n322), .ZN(n259) );
  NAND3_X1 U114 ( .A1(n354), .A2(n353), .A3(n352), .ZN(n356) );
  AOI21_X1 U115 ( .B1(\U4/DATA2_0 ), .B2(\U7/DATA1_0 ), .A(n328), .ZN(n327) );
  NAND2_X1 U116 ( .A1(n229), .A2(n394), .ZN(n395) );
  XOR2_X1 U117 ( .A(n367), .B(n366), .Z(n369) );
  XOR2_X1 U118 ( .A(n377), .B(n376), .Z(n378) );
  XOR2_X1 U119 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U120 ( .A1(n343), .A2(n342), .ZN(n346) );
  INV_X4 U121 ( .A(\U4/DATA2_18 ), .ZN(n392) );
  INV_X4 U122 ( .A(\U7/DATA1_18 ), .ZN(n271) );
  NAND2_X2 U123 ( .A1(n392), .A2(n271), .ZN(n309) );
  INV_X4 U124 ( .A(\U4/DATA2_16 ), .ZN(n273) );
  INV_X4 U125 ( .A(\U7/DATA1_16 ), .ZN(n272) );
  NAND2_X2 U126 ( .A1(n273), .A2(n272), .ZN(n306) );
  INV_X4 U127 ( .A(\U4/DATA2_15 ), .ZN(n275) );
  INV_X4 U128 ( .A(\U7/DATA1_15 ), .ZN(n274) );
  INV_X4 U129 ( .A(\U4/DATA2_14 ), .ZN(n277) );
  INV_X4 U130 ( .A(\U7/DATA1_14 ), .ZN(n276) );
  NAND2_X2 U131 ( .A1(n277), .A2(n276), .ZN(n305) );
  INV_X4 U132 ( .A(\U4/DATA2_13 ), .ZN(n279) );
  INV_X4 U133 ( .A(\U7/DATA1_13 ), .ZN(n278) );
  NAND2_X2 U134 ( .A1(n279), .A2(n278), .ZN(n303) );
  INV_X4 U135 ( .A(\U4/DATA2_12 ), .ZN(n281) );
  INV_X4 U136 ( .A(\U7/DATA1_12 ), .ZN(n280) );
  INV_X4 U137 ( .A(\U4/DATA2_11 ), .ZN(n283) );
  INV_X4 U138 ( .A(\U7/DATA1_11 ), .ZN(n282) );
  NAND2_X2 U139 ( .A1(n283), .A2(n282), .ZN(n302) );
  INV_X4 U140 ( .A(\U4/DATA2_10 ), .ZN(n285) );
  INV_X4 U141 ( .A(\U7/DATA1_10 ), .ZN(n284) );
  NAND2_X2 U142 ( .A1(n285), .A2(n284), .ZN(n300) );
  INV_X4 U143 ( .A(\U4/DATA2_9 ), .ZN(n287) );
  INV_X4 U144 ( .A(\U7/DATA1_9 ), .ZN(n286) );
  NAND2_X2 U145 ( .A1(n287), .A2(n286), .ZN(n298) );
  INV_X4 U146 ( .A(\U7/DATA1_8 ), .ZN(n288) );
  INV_X4 U147 ( .A(\U4/DATA2_7 ), .ZN(n364) );
  INV_X4 U148 ( .A(\U7/DATA1_7 ), .ZN(n407) );
  NAND2_X2 U149 ( .A1(n364), .A2(n407), .ZN(n293) );
  INV_X4 U150 ( .A(\U4/DATA2_4 ), .ZN(n344) );
  INV_X4 U151 ( .A(\U7/DATA1_4 ), .ZN(n404) );
  NAND2_X2 U152 ( .A1(n344), .A2(n404), .ZN(n352) );
  INV_X4 U153 ( .A(\U4/DATA2_5 ), .ZN(n350) );
  INV_X4 U154 ( .A(\U7/DATA1_5 ), .ZN(n405) );
  NAND2_X2 U155 ( .A1(n350), .A2(n405), .ZN(n354) );
  NAND2_X2 U156 ( .A1(\U4/DATA2_4 ), .A2(\U7/DATA1_4 ), .ZN(n348) );
  INV_X4 U157 ( .A(\U4/DATA2_1 ), .ZN(n329) );
  NAND2_X2 U158 ( .A1(n329), .A2(n402), .ZN(n289) );
  NAND2_X2 U159 ( .A1(n326), .A2(n401), .ZN(n325) );
  NAND2_X2 U160 ( .A1(n289), .A2(n325), .ZN(n331) );
  NAND2_X2 U161 ( .A1(\U4/DATA2_1 ), .A2(\U7/DATA1_1 ), .ZN(n332) );
  NAND2_X2 U162 ( .A1(\U4/DATA2_2 ), .A2(\U7/DATA1_2 ), .ZN(n338) );
  NAND2_X2 U163 ( .A1(n332), .A2(n338), .ZN(n290) );
  NAND3_X2 U164 ( .A1(n342), .A2(n348), .A3(n343), .ZN(n353) );
  NAND4_X2 U165 ( .A1(n293), .A2(n352), .A3(n354), .A4(n353), .ZN(n295) );
  NAND2_X2 U166 ( .A1(\U4/DATA2_5 ), .A2(\U7/DATA1_5 ), .ZN(n355) );
  NAND2_X2 U167 ( .A1(\U4/DATA2_6 ), .A2(\U7/DATA1_6 ), .ZN(n362) );
  NAND2_X2 U168 ( .A1(n355), .A2(n362), .ZN(n292) );
  NAND2_X2 U169 ( .A1(n293), .A2(n292), .ZN(n294) );
  INV_X4 U170 ( .A(\U4/DATA2_6 ), .ZN(n357) );
  INV_X4 U171 ( .A(\U7/DATA1_6 ), .ZN(n406) );
  NAND2_X2 U172 ( .A1(n357), .A2(n406), .ZN(n360) );
  NOR2_X2 U173 ( .A1(n407), .A2(n364), .ZN(n296) );
  AOI21_X4 U174 ( .B1(n297), .B2(n360), .A(n296), .ZN(n367) );
  AOI22_X4 U175 ( .A1(n237), .A2(n298), .B1(\U4/DATA2_9 ), .B2(\U7/DATA1_9 ), 
        .ZN(n372) );
  INV_X4 U176 ( .A(n372), .ZN(n299) );
  AOI22_X4 U177 ( .A1(n299), .A2(n300), .B1(\U4/DATA2_10 ), .B2(\U7/DATA1_10 ), 
        .ZN(n374) );
  INV_X4 U178 ( .A(n374), .ZN(n301) );
  AOI22_X4 U179 ( .A1(n301), .A2(n302), .B1(\U4/DATA2_11 ), .B2(\U7/DATA1_11 ), 
        .ZN(n377) );
  INV_X4 U180 ( .A(n381), .ZN(n304) );
  AOI22_X4 U181 ( .A1(n305), .A2(n304), .B1(\U7/DATA1_14 ), .B2(\U4/DATA2_14 ), 
        .ZN(n383) );
  AOI22_X4 U182 ( .A1(n306), .A2(n233), .B1(\U7/DATA1_16 ), .B2(\U4/DATA2_16 ), 
        .ZN(n388) );
  NOR2_X2 U183 ( .A1(\U7/DATA1_17 ), .A2(\U4/DATA2_17 ), .ZN(n308) );
  NAND2_X2 U184 ( .A1(\U7/DATA1_17 ), .A2(\U4/DATA2_17 ), .ZN(n307) );
  INV_X4 U185 ( .A(\U4/DATA2_19 ), .ZN(n398) );
  INV_X4 U186 ( .A(\U7/DATA1_19 ), .ZN(n310) );
  NAND2_X2 U187 ( .A1(n398), .A2(n310), .ZN(n319) );
  NAND2_X2 U188 ( .A1(\U7/DATA1_18 ), .A2(\U4/DATA2_18 ), .ZN(n394) );
  NAND2_X2 U189 ( .A1(\U7/DATA1_19 ), .A2(\U4/DATA2_19 ), .ZN(n312) );
  NAND2_X2 U190 ( .A1(divided[27]), .A2(n312), .ZN(n320) );
  INV_X4 U191 ( .A(n320), .ZN(n311) );
  INV_X4 U192 ( .A(n312), .ZN(n314) );
  INV_X4 U193 ( .A(divided[27]), .ZN(n313) );
  NAND2_X2 U194 ( .A1(n314), .A2(n313), .ZN(n315) );
  NAND3_X2 U195 ( .A1(n317), .A2(n316), .A3(n315), .ZN(n323) );
  INV_X4 U196 ( .A(n394), .ZN(n318) );
  NAND2_X2 U197 ( .A1(n318), .A2(n319), .ZN(n321) );
  OAI22_X2 U198 ( .A1(divided[27]), .A2(n321), .B1(n320), .B2(n319), .ZN(n322)
         );
  AND2_X1 U199 ( .A1(\U6/DATA1_6 ), .A2(n264), .ZN(\U6/Z_6 ) );
  OAI22_X2 U200 ( .A1(n327), .A2(n260), .B1(n262), .B2(n326), .ZN(n426) );
  OAI22_X2 U201 ( .A1(n330), .A2(n257), .B1(n329), .B2(n397), .ZN(n427) );
  OAI22_X2 U202 ( .A1(n334), .A2(n260), .B1(n333), .B2(n262), .ZN(n428) );
  NAND2_X2 U203 ( .A1(n336), .A2(n335), .ZN(n337) );
  XNOR2_X2 U204 ( .A(n340), .B(n339), .ZN(n341) );
  OAI22_X2 U205 ( .A1(n341), .A2(n257), .B1(n263), .B2(n254), .ZN(n409) );
  OAI22_X2 U206 ( .A1(n345), .A2(n399), .B1(n344), .B2(n263), .ZN(n410) );
  NAND2_X2 U207 ( .A1(n352), .A2(n346), .ZN(n347) );
  NAND2_X2 U208 ( .A1(n348), .A2(n347), .ZN(n349) );
  OAI22_X2 U209 ( .A1(n351), .A2(n260), .B1(n350), .B2(n397), .ZN(n411) );
  NAND2_X2 U210 ( .A1(n356), .A2(n355), .ZN(n359) );
  OAI22_X2 U211 ( .A1(n358), .A2(n257), .B1(n357), .B2(n262), .ZN(n412) );
  NAND2_X2 U212 ( .A1(n360), .A2(n359), .ZN(n361) );
  NAND2_X2 U213 ( .A1(n362), .A2(n361), .ZN(n363) );
  OAI22_X2 U214 ( .A1(n365), .A2(n399), .B1(n364), .B2(n263), .ZN(n413) );
  XOR2_X2 U215 ( .A(\U7/DATA1_8 ), .B(\U4/DATA2_8 ), .Z(n366) );
  INV_X4 U216 ( .A(\U4/DATA2_8 ), .ZN(n368) );
  OAI22_X2 U217 ( .A1(n369), .A2(n260), .B1(n368), .B2(n397), .ZN(n414) );
  OAI22_X2 U218 ( .A1(n371), .A2(n261), .B1(n287), .B2(n262), .ZN(n415) );
  OAI22_X2 U219 ( .A1(n373), .A2(n399), .B1(n285), .B2(n263), .ZN(n416) );
  OAI22_X2 U220 ( .A1(n375), .A2(n260), .B1(n283), .B2(n397), .ZN(n417) );
  XOR2_X2 U221 ( .A(\U7/DATA1_12 ), .B(\U4/DATA2_12 ), .Z(n376) );
  OAI22_X2 U222 ( .A1(n378), .A2(n261), .B1(n281), .B2(n262), .ZN(n418) );
  OAI22_X2 U223 ( .A1(n380), .A2(n399), .B1(n279), .B2(n263), .ZN(n419) );
  OAI22_X2 U224 ( .A1(n382), .A2(n260), .B1(n277), .B2(n397), .ZN(n420) );
  OAI22_X2 U225 ( .A1(n384), .A2(n261), .B1(n275), .B2(n262), .ZN(n421) );
  OAI22_X2 U226 ( .A1(n386), .A2(n399), .B1(n273), .B2(n263), .ZN(n422) );
  XOR2_X2 U227 ( .A(\U7/DATA1_17 ), .B(\U4/DATA2_17 ), .Z(n387) );
  INV_X4 U228 ( .A(\U4/DATA2_17 ), .ZN(n389) );
  OAI22_X2 U229 ( .A1(n390), .A2(n260), .B1(n389), .B2(n397), .ZN(n423) );
  OAI22_X2 U230 ( .A1(n393), .A2(n261), .B1(n392), .B2(n262), .ZN(n424) );
  XOR2_X2 U231 ( .A(\U7/DATA1_19 ), .B(\U4/DATA2_19 ), .Z(n396) );
  XNOR2_X2 U232 ( .A(n396), .B(n395), .ZN(n400) );
  OAI22_X2 U233 ( .A1(n400), .A2(n399), .B1(n398), .B2(n263), .ZN(n425) );
  NOR2_X2 U234 ( .A1(n265), .A2(n403), .ZN(\U7/Z_2 ) );
  NOR2_X2 U235 ( .A1(n265), .A2(n255), .ZN(\U7/Z_3 ) );
  NOR2_X2 U236 ( .A1(n265), .A2(n404), .ZN(\U7/Z_4 ) );
  NOR2_X2 U237 ( .A1(n265), .A2(n405), .ZN(\U7/Z_5 ) );
  NOR2_X2 U238 ( .A1(n265), .A2(n406), .ZN(\U7/Z_6 ) );
  NOR2_X2 U239 ( .A1(n265), .A2(n407), .ZN(\U7/Z_7 ) );
  NOR2_X2 U240 ( .A1(n265), .A2(n288), .ZN(\U7/Z_8 ) );
  NOR2_X2 U241 ( .A1(n265), .A2(n286), .ZN(\U7/Z_9 ) );
  NOR2_X2 U242 ( .A1(n265), .A2(n284), .ZN(\U7/Z_10 ) );
  NOR2_X2 U243 ( .A1(n282), .A2(n265), .ZN(\U7/Z_11 ) );
endmodule


module end_pipe_stage ( clock, reset_n, start, divided, divisor, q_in, 
        start_out, q_out );
  input [27:0] divided;
  input [19:0] divisor;
  input [7:0] q_in;
  output [7:0] q_out;
  input clock, reset_n, start;
  output start_out;
  wire   \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 , \U4/Z_7 ,
         \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 , \U4/DATA1_4 , \U4/DATA1_5 ,
         \U4/DATA1_6 , \U4/DATA1_7 , \stage_add/B[0] , \stage_add/B[1] ,
         \stage_add/B[2] , \stage_add/B[3] , \stage_add/B[4] ,
         \stage_add/B[5] , \stage_add/B[6] , \stage_add/B[7] ,
         \stage_add/B[8] , \stage_add/B[9] , \stage_add/B[10] ,
         \stage_add/B[11] , \stage_add/B[12] , \stage_add/B[13] ,
         \stage_add/B[14] , \stage_add/B[15] , \stage_add/B[16] ,
         \stage_add/B[17] , \stage_add/B[18] , \stage_add/B[19] ,
         \stage_add/A[0] , \stage_add/A[1] , \stage_add/A[2] ,
         \stage_add/A[3] , \stage_add/A[4] , \stage_add/A[5] ,
         \stage_add/A[6] , \stage_add/A[7] , \stage_add/A[8] ,
         \stage_add/A[9] , \stage_add/A[10] , \stage_add/A[11] ,
         \stage_add/A[12] , \stage_add/A[13] , \stage_add/A[14] ,
         \stage_add/A[15] , \stage_add/A[16] , \stage_add/A[17] ,
         \stage_add/A[18] , \stage_add/A[19] , n2, n105, n106, n107, n108,
         n109, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192;
  assign \U4/DATA1_1  = q_in[0];
  assign \U4/DATA1_2  = q_in[1];
  assign \U4/DATA1_3  = q_in[2];
  assign \U4/DATA1_4  = q_in[3];
  assign \U4/DATA1_5  = q_in[4];
  assign \U4/DATA1_6  = q_in[5];
  assign \U4/DATA1_7  = q_in[6];
  assign \stage_add/B[0]  = divisor[0];
  assign \stage_add/B[1]  = divisor[1];
  assign \stage_add/B[2]  = divisor[2];
  assign \stage_add/B[3]  = divisor[3];
  assign \stage_add/B[4]  = divisor[4];
  assign \stage_add/B[5]  = divisor[5];
  assign \stage_add/B[6]  = divisor[6];
  assign \stage_add/B[7]  = divisor[7];
  assign \stage_add/B[8]  = divisor[8];
  assign \stage_add/B[9]  = divisor[9];
  assign \stage_add/B[10]  = divisor[10];
  assign \stage_add/B[11]  = divisor[11];
  assign \stage_add/B[12]  = divisor[12];
  assign \stage_add/B[13]  = divisor[13];
  assign \stage_add/B[14]  = divisor[14];
  assign \stage_add/B[15]  = divisor[15];
  assign \stage_add/B[16]  = divisor[16];
  assign \stage_add/B[17]  = divisor[17];
  assign \stage_add/B[18]  = divisor[18];
  assign \stage_add/B[19]  = divisor[19];
  assign \stage_add/A[0]  = divided[7];
  assign \stage_add/A[1]  = divided[8];
  assign \stage_add/A[2]  = divided[9];
  assign \stage_add/A[3]  = divided[10];
  assign \stage_add/A[4]  = divided[11];
  assign \stage_add/A[5]  = divided[12];
  assign \stage_add/A[6]  = divided[13];
  assign \stage_add/A[7]  = divided[14];
  assign \stage_add/A[8]  = divided[15];
  assign \stage_add/A[9]  = divided[16];
  assign \stage_add/A[10]  = divided[17];
  assign \stage_add/A[11]  = divided[18];
  assign \stage_add/A[12]  = divided[19];
  assign \stage_add/A[13]  = divided[20];
  assign \stage_add/A[14]  = divided[21];
  assign \stage_add/A[15]  = divided[22];
  assign \stage_add/A[16]  = divided[23];
  assign \stage_add/A[17]  = divided[24];
  assign \stage_add/A[18]  = divided[25];
  assign \stage_add/A[19]  = divided[26];

  AND2_X1 U5 ( .A1(start), .A2(\U4/DATA1_7 ), .ZN(\U4/Z_7 ) );
  AND2_X1 U6 ( .A1(\U4/DATA1_6 ), .A2(start), .ZN(\U4/Z_6 ) );
  AND2_X1 U7 ( .A1(\U4/DATA1_5 ), .A2(start), .ZN(\U4/Z_5 ) );
  AND2_X1 U8 ( .A1(\U4/DATA1_4 ), .A2(start), .ZN(\U4/Z_4 ) );
  AND2_X1 U9 ( .A1(\U4/DATA1_3 ), .A2(start), .ZN(\U4/Z_3 ) );
  AND2_X1 U10 ( .A1(\U4/DATA1_2 ), .A2(start), .ZN(\U4/Z_2 ) );
  AND2_X1 U11 ( .A1(\U4/DATA1_1 ), .A2(start), .ZN(\U4/Z_1 ) );
  SDFFR_X1 \q_out_reg[0]  ( .D(start), .SI(1'b0), .SE(n2), .CK(clock), .RN(
        n121), .Q(q_out[0]) );
  DFFR_X2 start_out_reg ( .D(start), .CK(clock), .RN(n121), .Q(start_out) );
  DFFR_X2 \q_out_reg[7]  ( .D(\U4/Z_7 ), .CK(clock), .RN(n121), .Q(q_out[7])
         );
  DFFR_X2 \q_out_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n121), .Q(q_out[6])
         );
  DFFR_X2 \q_out_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n121), .Q(q_out[5])
         );
  DFFR_X2 \q_out_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(n121), .Q(q_out[4])
         );
  DFFR_X2 \q_out_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n121), .Q(q_out[3])
         );
  DFFR_X2 \q_out_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .RN(n121), .Q(q_out[2])
         );
  DFFR_X2 \q_out_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .RN(n121), .Q(q_out[1])
         );
  AOI22_X2 U4 ( .A1(n106), .A2(n109), .B1(n107), .B2(n108), .ZN(n105) );
  INV_X32 U12 ( .A(n179), .ZN(n106) );
  INV_X32 U13 ( .A(\stage_add/B[17] ), .ZN(n107) );
  INV_X32 U14 ( .A(\stage_add/A[17] ), .ZN(n108) );
  NAND2_X2 U15 ( .A1(\stage_add/A[16] ), .A2(\stage_add/B[16] ), .ZN(n109) );
  OAI21_X2 U16 ( .B1(n147), .B2(n112), .A(n146), .ZN(n150) );
  OAI211_X2 U17 ( .C1(n119), .C2(n120), .A(n131), .B(n132), .ZN(n118) );
  AND2_X4 U18 ( .A1(\stage_add/A[4] ), .A2(\stage_add/B[4] ), .ZN(n111) );
  AND2_X4 U19 ( .A1(\stage_add/A[6] ), .A2(\stage_add/B[6] ), .ZN(n112) );
  AND2_X4 U20 ( .A1(\stage_add/A[8] ), .A2(\stage_add/B[8] ), .ZN(n113) );
  AND2_X4 U21 ( .A1(\stage_add/A[10] ), .A2(\stage_add/B[10] ), .ZN(n114) );
  AND2_X4 U22 ( .A1(\stage_add/A[12] ), .A2(\stage_add/B[12] ), .ZN(n115) );
  AND2_X4 U23 ( .A1(\stage_add/A[14] ), .A2(\stage_add/B[14] ), .ZN(n116) );
  AND2_X4 U24 ( .A1(\stage_add/B[18] ), .A2(\stage_add/A[18] ), .ZN(n117) );
  OAI21_X4 U25 ( .B1(n140), .B2(n111), .A(n139), .ZN(n143) );
  OAI21_X4 U26 ( .B1(n105), .B2(n185), .A(n184), .ZN(n190) );
  INV_X1 U27 ( .A(n133), .ZN(n120) );
  INV_X4 U28 ( .A(n118), .ZN(n136) );
  INV_X4 U29 ( .A(n134), .ZN(n119) );
  NAND3_X2 U30 ( .A1(\stage_add/B[2] ), .A2(\stage_add/A[2] ), .A3(n133), .ZN(
        n132) );
  NAND2_X1 U31 ( .A1(\stage_add/B[3] ), .A2(\stage_add/A[3] ), .ZN(n131) );
  OR2_X2 U32 ( .A1(\stage_add/A[3] ), .A2(\stage_add/B[3] ), .ZN(n133) );
  INV_X4 U33 ( .A(n122), .ZN(n121) );
  INV_X4 U34 ( .A(reset_n), .ZN(n122) );
  AOI21_X2 U35 ( .B1(n130), .B2(n129), .A(n128), .ZN(n134) );
  AOI21_X2 U36 ( .B1(n143), .B2(n142), .A(n141), .ZN(n147) );
  OAI21_X2 U37 ( .B1(n154), .B2(n113), .A(n153), .ZN(n157) );
  AOI21_X2 U38 ( .B1(n150), .B2(n149), .A(n148), .ZN(n154) );
  OAI21_X2 U39 ( .B1(n161), .B2(n114), .A(n160), .ZN(n164) );
  AOI21_X2 U40 ( .B1(n157), .B2(n156), .A(n155), .ZN(n161) );
  OAI21_X2 U41 ( .B1(n168), .B2(n115), .A(n167), .ZN(n171) );
  AOI21_X2 U42 ( .B1(n164), .B2(n163), .A(n162), .ZN(n168) );
  OAI21_X2 U43 ( .B1(n175), .B2(n116), .A(n174), .ZN(n178) );
  AOI21_X2 U44 ( .B1(n171), .B2(n170), .A(n169), .ZN(n175) );
  AOI21_X2 U45 ( .B1(n178), .B2(n177), .A(n176), .ZN(n179) );
  NAND2_X2 U46 ( .A1(\stage_add/B[19] ), .A2(\stage_add/A[19] ), .ZN(n127) );
  NAND2_X2 U47 ( .A1(divided[27]), .A2(n127), .ZN(n187) );
  INV_X4 U48 ( .A(\stage_add/A[19] ), .ZN(n124) );
  INV_X4 U49 ( .A(\stage_add/B[19] ), .ZN(n123) );
  NAND2_X2 U50 ( .A1(n124), .A2(n123), .ZN(n186) );
  INV_X4 U51 ( .A(divided[27]), .ZN(n125) );
  NAND3_X2 U52 ( .A1(n117), .A2(n186), .A3(n125), .ZN(n126) );
  OAI221_X2 U53 ( .B1(n187), .B2(n186), .C1(divided[27]), .C2(n127), .A(n126), 
        .ZN(n192) );
  NAND2_X2 U54 ( .A1(\stage_add/B[1] ), .A2(\stage_add/A[1] ), .ZN(n130) );
  OAI22_X2 U55 ( .A1(\stage_add/B[1] ), .A2(\stage_add/A[1] ), .B1(
        \stage_add/B[0] ), .B2(\stage_add/A[0] ), .ZN(n129) );
  NOR2_X2 U56 ( .A1(\stage_add/B[2] ), .A2(\stage_add/A[2] ), .ZN(n128) );
  NOR2_X2 U57 ( .A1(\stage_add/B[4] ), .A2(\stage_add/A[4] ), .ZN(n135) );
  NOR2_X2 U58 ( .A1(n136), .A2(n135), .ZN(n140) );
  INV_X4 U59 ( .A(\stage_add/A[5] ), .ZN(n138) );
  INV_X4 U60 ( .A(\stage_add/B[5] ), .ZN(n137) );
  NAND2_X2 U61 ( .A1(n138), .A2(n137), .ZN(n139) );
  NAND2_X2 U62 ( .A1(\stage_add/B[5] ), .A2(\stage_add/A[5] ), .ZN(n142) );
  NOR2_X2 U63 ( .A1(\stage_add/B[6] ), .A2(\stage_add/A[6] ), .ZN(n141) );
  INV_X4 U64 ( .A(\stage_add/A[7] ), .ZN(n145) );
  INV_X4 U65 ( .A(\stage_add/B[7] ), .ZN(n144) );
  NAND2_X2 U66 ( .A1(n145), .A2(n144), .ZN(n146) );
  NAND2_X2 U67 ( .A1(\stage_add/B[7] ), .A2(\stage_add/A[7] ), .ZN(n149) );
  NOR2_X2 U68 ( .A1(\stage_add/B[8] ), .A2(\stage_add/A[8] ), .ZN(n148) );
  INV_X4 U69 ( .A(\stage_add/A[9] ), .ZN(n152) );
  INV_X4 U70 ( .A(\stage_add/B[9] ), .ZN(n151) );
  NAND2_X2 U71 ( .A1(n152), .A2(n151), .ZN(n153) );
  NAND2_X2 U72 ( .A1(\stage_add/B[9] ), .A2(\stage_add/A[9] ), .ZN(n156) );
  NOR2_X2 U73 ( .A1(\stage_add/B[10] ), .A2(\stage_add/A[10] ), .ZN(n155) );
  INV_X4 U74 ( .A(\stage_add/A[11] ), .ZN(n159) );
  INV_X4 U75 ( .A(\stage_add/B[11] ), .ZN(n158) );
  NAND2_X2 U76 ( .A1(n159), .A2(n158), .ZN(n160) );
  NAND2_X2 U77 ( .A1(\stage_add/B[11] ), .A2(\stage_add/A[11] ), .ZN(n163) );
  NOR2_X2 U78 ( .A1(\stage_add/B[12] ), .A2(\stage_add/A[12] ), .ZN(n162) );
  INV_X4 U79 ( .A(\stage_add/A[13] ), .ZN(n166) );
  INV_X4 U80 ( .A(\stage_add/B[13] ), .ZN(n165) );
  NAND2_X2 U81 ( .A1(n166), .A2(n165), .ZN(n167) );
  NAND2_X2 U82 ( .A1(\stage_add/B[13] ), .A2(\stage_add/A[13] ), .ZN(n170) );
  NOR2_X2 U83 ( .A1(\stage_add/B[14] ), .A2(\stage_add/A[14] ), .ZN(n169) );
  INV_X4 U84 ( .A(\stage_add/A[15] ), .ZN(n173) );
  INV_X4 U85 ( .A(\stage_add/B[15] ), .ZN(n172) );
  NAND2_X2 U86 ( .A1(n173), .A2(n172), .ZN(n174) );
  NAND2_X2 U87 ( .A1(\stage_add/B[15] ), .A2(\stage_add/A[15] ), .ZN(n177) );
  NOR2_X2 U88 ( .A1(\stage_add/B[16] ), .A2(\stage_add/A[16] ), .ZN(n176) );
  INV_X4 U89 ( .A(\stage_add/A[17] ), .ZN(n181) );
  INV_X4 U90 ( .A(\stage_add/B[17] ), .ZN(n180) );
  NOR2_X2 U91 ( .A1(n181), .A2(n180), .ZN(n185) );
  INV_X4 U92 ( .A(\stage_add/A[18] ), .ZN(n183) );
  INV_X4 U93 ( .A(\stage_add/B[18] ), .ZN(n182) );
  NAND2_X2 U94 ( .A1(n183), .A2(n182), .ZN(n184) );
  INV_X4 U95 ( .A(n186), .ZN(n189) );
  INV_X4 U96 ( .A(n190), .ZN(n188) );
  OAI33_X1 U97 ( .A1(n190), .A2(divided[27]), .A3(n189), .B1(n188), .B2(n117), 
        .B3(n187), .ZN(n191) );
  NOR2_X2 U98 ( .A1(n191), .A2(n192), .ZN(n2) );
endmodule


module pipeline_divider ( clock, reset_n, start, divided, divisor, q, StartOut
 );
  input [27:0] divided;
  input [19:0] divisor;
  output [7:0] q;
  input clock, reset_n, start;
  output StartOut;
  wire   start1, start2, start3, start4, start5, start6, start7, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22;
  wire   [19:0] divisor1;
  wire   [27:0] result1;
  wire   [7:0] q0;
  wire   [19:0] divisor2;
  wire   [27:0] result2;
  wire   [7:0] q1;
  wire   [19:0] divisor3;
  wire   [27:0] result3;
  wire   [7:0] q2;
  wire   [19:0] divisor4;
  wire   [27:0] result4;
  wire   [7:0] q3;
  wire   [19:0] divisor5;
  wire   [27:0] result5;
  wire   [7:0] q4;
  wire   [19:0] divisor6;
  wire   [27:0] result6;
  wire   [7:0] q5;
  wire   [19:0] divisor7;
  wire   [27:0] result7;
  wire   [7:0] q6;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  divider_pipe_stage_1 stage0 ( .clock(clock), .reset_n(n21), .start(start), 
        .divided(divided), .divisor({n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
        n11, n12, n13, n14, n15, n16, n17, n18, n19, n20}), .q_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .start_out(start1), 
        .divisor_out(divisor1), .result({result1[27:1], 
        SYNOPSYS_UNCONNECTED__0}), .q_out(q0) );
  divider_pipe_stage_6 stage1 ( .clock(clock), .reset_n(n21), .start(start1), 
        .divided({result1[27:1], 1'b0}), .divisor(divisor1), .q_in(q0), 
        .start_out(start2), .divisor_out(divisor2), .result({result2[27:1], 
        SYNOPSYS_UNCONNECTED__1}), .q_out(q1) );
  divider_pipe_stage_5 stage2 ( .clock(clock), .reset_n(n21), .start(start2), 
        .divided({result2[27:1], 1'b0}), .divisor(divisor2), .q_in(q1), 
        .start_out(start3), .divisor_out(divisor3), .result({result3[27:1], 
        SYNOPSYS_UNCONNECTED__2}), .q_out(q2) );
  divider_pipe_stage_4 stage3 ( .clock(clock), .reset_n(n21), .start(start3), 
        .divided({result3[27:1], 1'b0}), .divisor(divisor3), .q_in(q2), 
        .start_out(start4), .divisor_out(divisor4), .result({result4[27:1], 
        SYNOPSYS_UNCONNECTED__3}), .q_out(q3) );
  divider_pipe_stage_3 stage4 ( .clock(clock), .reset_n(n21), .start(start4), 
        .divided({result4[27:1], 1'b0}), .divisor(divisor4), .q_in(q3), 
        .start_out(start5), .divisor_out(divisor5), .result({result5[27:1], 
        SYNOPSYS_UNCONNECTED__4}), .q_out(q4) );
  divider_pipe_stage_2 stage5 ( .clock(clock), .reset_n(n21), .start(start5), 
        .divided({result5[27:1], 1'b0}), .divisor(divisor5), .q_in(q4), 
        .start_out(start6), .divisor_out(divisor6), .result({result6[27:1], 
        SYNOPSYS_UNCONNECTED__5}), .q_out(q5) );
  divider_pipe_stage_0 stage6 ( .clock(clock), .reset_n(n21), .start(start6), 
        .divided({result6[27:1], 1'b0}), .divisor(divisor6), .q_in(q5), 
        .start_out(start7), .divisor_out(divisor7), .result({result7[27:1], 
        SYNOPSYS_UNCONNECTED__6}), .q_out(q6) );
  end_pipe_stage stage7 ( .clock(clock), .reset_n(n21), .start(start7), 
        .divided({result7[27:1], 1'b0}), .divisor(divisor7), .q_in(q6), 
        .start_out(StartOut), .q_out(q) );
  INV_X2 U2 ( .A(divisor[15]), .ZN(n5) );
  INV_X4 U3 ( .A(n22), .ZN(n21) );
  INV_X4 U4 ( .A(reset_n), .ZN(n22) );
  INV_X4 U5 ( .A(divisor[0]), .ZN(n20) );
  INV_X4 U6 ( .A(divisor[1]), .ZN(n19) );
  INV_X4 U7 ( .A(divisor[2]), .ZN(n18) );
  INV_X4 U8 ( .A(divisor[3]), .ZN(n17) );
  INV_X4 U9 ( .A(divisor[4]), .ZN(n16) );
  INV_X4 U10 ( .A(divisor[5]), .ZN(n15) );
  INV_X4 U11 ( .A(divisor[6]), .ZN(n14) );
  INV_X4 U12 ( .A(divisor[7]), .ZN(n13) );
  INV_X4 U13 ( .A(divisor[8]), .ZN(n12) );
  INV_X4 U14 ( .A(divisor[9]), .ZN(n11) );
  INV_X4 U15 ( .A(divisor[10]), .ZN(n10) );
  INV_X4 U16 ( .A(divisor[11]), .ZN(n9) );
  INV_X4 U17 ( .A(divisor[12]), .ZN(n8) );
  INV_X4 U18 ( .A(divisor[13]), .ZN(n7) );
  INV_X4 U19 ( .A(divisor[14]), .ZN(n6) );
  INV_X4 U20 ( .A(divisor[16]), .ZN(n4) );
  INV_X4 U21 ( .A(divisor[17]), .ZN(n3) );
  INV_X4 U22 ( .A(divisor[18]), .ZN(n2) );
  INV_X4 U23 ( .A(divisor[19]), .ZN(n1) );
endmodule


module Output_Result ( clock, reset_n, DataIn, StartIn, Divisor, StartOut, 
        DataOut );
  input [27:0] DataIn;
  input [19:0] Divisor;
  output [7:0] DataOut;
  input clock, reset_n, StartIn;
  output StartOut;


  pipeline_divider divider ( .clock(clock), .reset_n(reset_n), .start(StartIn), 
        .divided(DataIn), .divisor(Divisor), .q(DataOut), .StartOut(StartOut)
         );
endmodule


module Output_Store ( clock, reset_n, StartIn, ResultIn, WriteBus, 
        WriteAddress, WriteEnable, output_base_offset );
  input [7:0] ResultIn;
  output [127:0] WriteBus;
  output [15:0] WriteAddress;
  input clock, reset_n, StartIn, output_base_offset;
  output WriteEnable;
  wire   \U8/DATA1_0 , \U8/DATA1_1 , \U8/DATA1_2 , \U8/DATA1_3 , \U8/DATA1_4 ,
         \U8/DATA1_5 , \U8/DATA1_6 , \U8/DATA1_7 , \U7/Z_0 , \U7/Z_1 ,
         \U7/Z_2 , \U7/Z_3 , \U6/Z_0 , \U5/DATA2_1 , \U5/DATA2_2 ,
         \U5/DATA2_3 , \U5/DATA2_4 , \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 ,
         \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 , \U4/DATA1_7 , \U4/DATA1_8 ,
         \U4/DATA1_9 , \U4/DATA1_10 , \U4/DATA1_11 , \U4/DATA1_12 ,
         \U4/DATA1_13 , \U4/DATA1_14 , \sub_63/carry[2] , \sub_63/carry[3] ,
         \sub_63/carry[4] , \sub_63/A[0] , \sub_63/A[1] , \sub_63/A[2] ,
         \sub_63/A[3] , \sub_63/A[4] , \add_55/carry[15] , \add_55/carry[12] ,
         \add_55/carry[11] , \add_55/carry[9] , \add_55/carry[8] ,
         \add_55/carry[7] , \add_55/carry[6] , \add_55/carry[5] ,
         \add_55/carry[3] , \add_55/carry[2] , \add_55/A[0] , \add_55/A[1] ,
         \add_55/A[2] , \add_55/A[3] , \add_55/A[4] , \add_55/A[5] ,
         \add_55/A[6] , \add_55/A[7] , \add_55/A[8] , \add_55/A[9] ,
         \add_55/A[10] , \add_55/A[11] , \add_55/A[12] , \add_55/A[13] ,
         \add_55/A[14] , \add_55/A[15] , n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n133, n135, n136, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571;
  assign \U8/DATA1_0  = ResultIn[0];
  assign \U8/DATA1_1  = ResultIn[1];
  assign \U8/DATA1_2  = ResultIn[2];
  assign \U8/DATA1_3  = ResultIn[3];
  assign \U8/DATA1_4  = ResultIn[4];
  assign \U8/DATA1_5  = ResultIn[5];
  assign \U8/DATA1_6  = ResultIn[6];
  assign \U8/DATA1_7  = ResultIn[7];

  HA_X1 \add_55/U1_1_1  ( .A(\add_55/A[1] ), .B(\add_55/A[0] ), .CO(
        \add_55/carry[2] ), .S(\U4/DATA1_1 ) );
  HA_X1 \add_55/U1_1_2  ( .A(\add_55/A[2] ), .B(\add_55/carry[2] ), .CO(
        \add_55/carry[3] ), .S(\U4/DATA1_2 ) );
  HA_X1 \add_55/U1_1_4  ( .A(\add_55/A[4] ), .B(n494), .CO(\add_55/carry[5] ), 
        .S(\U4/DATA1_4 ) );
  HA_X1 \add_55/U1_1_5  ( .A(\add_55/A[5] ), .B(\add_55/carry[5] ), .CO(
        \add_55/carry[6] ), .S(\U4/DATA1_5 ) );
  HA_X1 \add_55/U1_1_6  ( .A(\add_55/A[6] ), .B(\add_55/carry[6] ), .CO(
        \add_55/carry[7] ), .S(\U4/DATA1_6 ) );
  HA_X1 \add_55/U1_1_7  ( .A(\add_55/A[7] ), .B(\add_55/carry[7] ), .CO(
        \add_55/carry[8] ), .S(\U4/DATA1_7 ) );
  HA_X1 \add_55/U1_1_8  ( .A(\add_55/A[8] ), .B(\add_55/carry[8] ), .CO(
        \add_55/carry[9] ), .S(\U4/DATA1_8 ) );
  HA_X1 \add_55/U1_1_10  ( .A(\add_55/A[10] ), .B(n493), .CO(
        \add_55/carry[11] ), .S(\U4/DATA1_10 ) );
  HA_X1 \add_55/U1_1_11  ( .A(\add_55/A[11] ), .B(\add_55/carry[11] ), .CO(
        \add_55/carry[12] ), .S(\U4/DATA1_11 ) );
  HA_X1 \add_55/U1_1_14  ( .A(\add_55/A[14] ), .B(n492), .CO(
        \add_55/carry[15] ), .S(\U4/DATA1_14 ) );
  XNOR2_X2 \sub_63/U1_A_1  ( .A(\sub_63/A[1] ), .B(\sub_63/A[0] ), .ZN(
        \U5/DATA2_1 ) );
  OR2_X1 \sub_63/U1_B_1  ( .A1(\sub_63/A[1] ), .A2(\sub_63/A[0] ), .ZN(
        \sub_63/carry[2] ) );
  XNOR2_X2 \sub_63/U1_A_2  ( .A(\sub_63/A[2] ), .B(\sub_63/carry[2] ), .ZN(
        \U5/DATA2_2 ) );
  OR2_X1 \sub_63/U1_B_2  ( .A1(\sub_63/A[2] ), .A2(\sub_63/carry[2] ), .ZN(
        \sub_63/carry[3] ) );
  XNOR2_X2 \sub_63/U1_A_3  ( .A(\sub_63/A[3] ), .B(\sub_63/carry[3] ), .ZN(
        \U5/DATA2_3 ) );
  OR2_X1 \sub_63/U1_B_3  ( .A1(\sub_63/A[3] ), .A2(\sub_63/carry[3] ), .ZN(
        \sub_63/carry[4] ) );
  XNOR2_X2 \sub_63/U1_A_4  ( .A(\sub_63/A[4] ), .B(\sub_63/carry[4] ), .ZN(
        \U5/DATA2_4 ) );
  DFFS_X2 \short_count_reg[0]  ( .D(\U7/Z_0 ), .CK(clock), .SN(n511), .Q(
        \sub_63/A[0] ), .QN(n66) );
  DFFS_X2 \short_count_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .SN(n511), .Q(
        \sub_63/A[1] ), .QN(n65) );
  DFFS_X2 \short_count_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .SN(n511), .Q(
        \sub_63/A[2] ), .QN(n64) );
  DFFS_X2 \short_count_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .SN(n511), .Q(
        \sub_63/A[3] ), .QN(n63) );
  SDFFR_X2 \short_count_reg[4]  ( .D(1'b0), .SI(n549), .SE(\U5/DATA2_4 ), .CK(
        clock), .RN(n511), .Q(\sub_63/A[4] ) );
  DFFR_X1 \next_WriteAddress_reg[3]  ( .D(n516), .CK(clock), .RN(n511), .Q(
        \add_55/A[3] ) );
  DFFR_X1 \next_WriteAddress_reg[4]  ( .D(n517), .CK(clock), .RN(n511), .Q(
        \add_55/A[4] ) );
  DFFR_X1 \next_WriteAddress_reg[5]  ( .D(n518), .CK(clock), .RN(n511), .Q(
        \add_55/A[5] ) );
  DFFR_X1 \next_WriteAddress_reg[6]  ( .D(n519), .CK(clock), .RN(n503), .Q(
        \add_55/A[6] ) );
  DFFR_X1 \next_WriteAddress_reg[7]  ( .D(n520), .CK(clock), .RN(n511), .Q(
        \add_55/A[7] ) );
  DFFR_X1 \next_WriteAddress_reg[8]  ( .D(n521), .CK(clock), .RN(n511), .Q(
        \add_55/A[8] ) );
  DFFR_X1 \next_WriteAddress_reg[9]  ( .D(n522), .CK(clock), .RN(n511), .Q(
        \add_55/A[9] ) );
  DFFR_X1 \next_WriteAddress_reg[10]  ( .D(n523), .CK(clock), .RN(n511), .Q(
        \add_55/A[10] ) );
  DFFR_X1 \next_WriteAddress_reg[11]  ( .D(n524), .CK(clock), .RN(n511), .Q(
        \add_55/A[11] ) );
  DFFR_X1 \next_WriteAddress_reg[12]  ( .D(n525), .CK(clock), .RN(n511), .Q(
        \add_55/A[12] ) );
  NAND3_X2 U5 ( .A1(n498), .A2(n130), .A3(\add_55/carry[15] ), .ZN(n133) );
  OAI22_X2 U23 ( .A1(n539), .A2(n151), .B1(n152), .B2(n129), .ZN(n362) );
  OAI22_X2 U24 ( .A1(n539), .A2(n153), .B1(n152), .B2(n128), .ZN(n363) );
  OAI22_X2 U25 ( .A1(n539), .A2(n154), .B1(n152), .B2(n127), .ZN(n364) );
  OAI22_X2 U26 ( .A1(n539), .A2(n155), .B1(n152), .B2(n126), .ZN(n365) );
  OAI22_X2 U27 ( .A1(n539), .A2(n156), .B1(n152), .B2(n125), .ZN(n366) );
  OAI22_X2 U28 ( .A1(n539), .A2(n157), .B1(n152), .B2(n124), .ZN(n367) );
  OAI22_X2 U29 ( .A1(n539), .A2(n158), .B1(n152), .B2(n123), .ZN(n368) );
  OAI22_X2 U30 ( .A1(n539), .A2(n159), .B1(n152), .B2(n122), .ZN(n369) );
  NAND2_X2 U31 ( .A1(n499), .A2(n160), .ZN(n152) );
  NAND4_X2 U32 ( .A1(n161), .A2(n162), .A3(n163), .A4(n164), .ZN(n160) );
  OAI22_X2 U33 ( .A1(n538), .A2(n151), .B1(n165), .B2(n121), .ZN(n370) );
  NAND2_X2 U34 ( .A1(n499), .A2(n166), .ZN(n165) );
  NAND3_X2 U35 ( .A1(n161), .A2(n167), .A3(n557), .ZN(n166) );
  OAI22_X2 U36 ( .A1(n153), .A2(n168), .B1(n534), .B2(n120), .ZN(n371) );
  NAND2_X2 U37 ( .A1(n169), .A2(n170), .ZN(n168) );
  NAND2_X2 U40 ( .A1(WriteBus[10]), .A2(n173), .ZN(n174) );
  NAND2_X2 U42 ( .A1(WriteBus[11]), .A2(n173), .ZN(n175) );
  NAND2_X2 U44 ( .A1(WriteBus[12]), .A2(n173), .ZN(n176) );
  NAND2_X2 U46 ( .A1(WriteBus[13]), .A2(n173), .ZN(n177) );
  NAND2_X2 U48 ( .A1(WriteBus[14]), .A2(n173), .ZN(n178) );
  NOR4_X2 U50 ( .A1(n566), .A2(n547), .A3(n180), .A4(n181), .ZN(n179) );
  NAND2_X2 U52 ( .A1(WriteBus[15]), .A2(n182), .ZN(n183) );
  NAND4_X2 U53 ( .A1(n540), .A2(n184), .A3(n527), .A4(n185), .ZN(n182) );
  NAND3_X2 U55 ( .A1(n189), .A2(n190), .A3(n191), .ZN(n186) );
  NAND2_X2 U58 ( .A1(WriteBus[16]), .A2(n195), .ZN(n196) );
  NAND2_X2 U60 ( .A1(WriteBus[17]), .A2(n195), .ZN(n197) );
  NAND2_X2 U62 ( .A1(WriteBus[18]), .A2(n195), .ZN(n198) );
  NAND2_X2 U64 ( .A1(WriteBus[19]), .A2(n195), .ZN(n199) );
  NAND2_X2 U66 ( .A1(WriteBus[20]), .A2(n195), .ZN(n200) );
  NAND2_X2 U68 ( .A1(WriteBus[21]), .A2(n195), .ZN(n201) );
  NOR3_X2 U70 ( .A1(n205), .A2(n570), .A3(n206), .ZN(n202) );
  NAND2_X2 U72 ( .A1(WriteBus[22]), .A2(n207), .ZN(n208) );
  NAND2_X2 U74 ( .A1(WriteBus[23]), .A2(n207), .ZN(n209) );
  NAND3_X2 U75 ( .A1(n210), .A2(n211), .A3(n204), .ZN(n207) );
  NAND2_X2 U77 ( .A1(WriteBus[24]), .A2(n212), .ZN(n213) );
  NAND2_X2 U79 ( .A1(WriteBus[25]), .A2(n212), .ZN(n214) );
  NAND2_X2 U81 ( .A1(WriteBus[26]), .A2(n212), .ZN(n215) );
  NAND2_X2 U83 ( .A1(WriteBus[27]), .A2(n212), .ZN(n216) );
  NAND2_X2 U85 ( .A1(WriteBus[28]), .A2(n212), .ZN(n217) );
  NOR3_X2 U87 ( .A1(n206), .A2(n564), .A3(n570), .ZN(n218) );
  OAI22_X2 U88 ( .A1(n537), .A2(n157), .B1(n219), .B2(n119), .ZN(n391) );
  OAI22_X2 U89 ( .A1(n537), .A2(n158), .B1(n219), .B2(n118), .ZN(n392) );
  OAI22_X2 U90 ( .A1(n537), .A2(n159), .B1(n219), .B2(n117), .ZN(n393) );
  NAND2_X2 U91 ( .A1(n499), .A2(n220), .ZN(n219) );
  NAND4_X2 U92 ( .A1(n555), .A2(n161), .A3(n163), .A4(n221), .ZN(n220) );
  OAI22_X2 U93 ( .A1(n536), .A2(n151), .B1(n222), .B2(n116), .ZN(n394) );
  OAI22_X2 U94 ( .A1(n536), .A2(n153), .B1(n222), .B2(n115), .ZN(n395) );
  OAI22_X2 U95 ( .A1(n536), .A2(n154), .B1(n222), .B2(n114), .ZN(n396) );
  OAI22_X2 U96 ( .A1(n536), .A2(n155), .B1(n222), .B2(n113), .ZN(n397) );
  OAI22_X2 U97 ( .A1(n536), .A2(n156), .B1(n222), .B2(n112), .ZN(n398) );
  OAI22_X2 U98 ( .A1(n536), .A2(n157), .B1(n222), .B2(n111), .ZN(n399) );
  OAI22_X2 U99 ( .A1(n536), .A2(n158), .B1(n222), .B2(n110), .ZN(n400) );
  OAI22_X2 U100 ( .A1(n536), .A2(n159), .B1(n222), .B2(n109), .ZN(n401) );
  NAND2_X2 U101 ( .A1(n499), .A2(n223), .ZN(n222) );
  NAND4_X2 U102 ( .A1(n557), .A2(n161), .A3(n224), .A4(n164), .ZN(n223) );
  NAND2_X2 U104 ( .A1(WriteBus[40]), .A2(n225), .ZN(n226) );
  NAND2_X2 U106 ( .A1(WriteBus[41]), .A2(n225), .ZN(n227) );
  AND3_X2 U108 ( .A1(n184), .A2(n229), .A3(n230), .ZN(n161) );
  OAI22_X2 U109 ( .A1(n154), .A2(n231), .B1(n533), .B2(n108), .ZN(n404) );
  OAI22_X2 U110 ( .A1(n155), .A2(n231), .B1(n533), .B2(n107), .ZN(n405) );
  OAI22_X2 U111 ( .A1(n156), .A2(n231), .B1(n533), .B2(n106), .ZN(n406) );
  OAI22_X2 U112 ( .A1(n157), .A2(n231), .B1(n533), .B2(n105), .ZN(n407) );
  OAI22_X2 U113 ( .A1(n158), .A2(n231), .B1(n533), .B2(n104), .ZN(n408) );
  OAI22_X2 U114 ( .A1(n159), .A2(n231), .B1(n533), .B2(n103), .ZN(n409) );
  NAND2_X2 U115 ( .A1(n169), .A2(n232), .ZN(n231) );
  NAND3_X2 U117 ( .A1(n234), .A2(n164), .A3(n557), .ZN(n228) );
  OAI22_X2 U118 ( .A1(n151), .A2(n235), .B1(n532), .B2(n102), .ZN(n410) );
  NAND3_X2 U119 ( .A1(n236), .A2(n237), .A3(n169), .ZN(n235) );
  NAND2_X2 U122 ( .A1(WriteBus[49]), .A2(n238), .ZN(n239) );
  NAND2_X2 U124 ( .A1(WriteBus[50]), .A2(n238), .ZN(n240) );
  NAND2_X2 U126 ( .A1(WriteBus[51]), .A2(n238), .ZN(n241) );
  NAND2_X2 U128 ( .A1(WriteBus[52]), .A2(n238), .ZN(n242) );
  NAND2_X2 U130 ( .A1(WriteBus[53]), .A2(n238), .ZN(n243) );
  NAND2_X2 U132 ( .A1(WriteBus[54]), .A2(n238), .ZN(n244) );
  NOR3_X2 U134 ( .A1(n247), .A2(n561), .A3(n172), .ZN(n245) );
  NAND2_X2 U136 ( .A1(WriteBus[55]), .A2(n248), .ZN(n249) );
  NAND3_X2 U137 ( .A1(n250), .A2(n251), .A3(n246), .ZN(n248) );
  NAND2_X2 U140 ( .A1(WriteBus[56]), .A2(n252), .ZN(n253) );
  NAND2_X2 U142 ( .A1(WriteBus[57]), .A2(n252), .ZN(n254) );
  NAND2_X2 U144 ( .A1(WriteBus[58]), .A2(n252), .ZN(n255) );
  NAND2_X2 U146 ( .A1(WriteBus[59]), .A2(n252), .ZN(n256) );
  NAND2_X2 U148 ( .A1(WriteBus[60]), .A2(n252), .ZN(n257) );
  NAND2_X2 U150 ( .A1(WriteBus[61]), .A2(n252), .ZN(n258) );
  NOR3_X2 U152 ( .A1(n261), .A2(n247), .A3(n262), .ZN(n259) );
  NAND3_X2 U153 ( .A1(n263), .A2(n565), .A3(n221), .ZN(n261) );
  OAI22_X2 U154 ( .A1(n158), .A2(n264), .B1(n529), .B2(n101), .ZN(n424) );
  OAI22_X2 U155 ( .A1(n159), .A2(n264), .B1(n529), .B2(n100), .ZN(n425) );
  NAND3_X2 U156 ( .A1(n230), .A2(n184), .A3(n265), .ZN(n264) );
  OAI22_X2 U157 ( .A1(n151), .A2(n266), .B1(n528), .B2(n99), .ZN(n426) );
  OAI22_X2 U158 ( .A1(n153), .A2(n266), .B1(n528), .B2(n98), .ZN(n427) );
  OAI22_X2 U159 ( .A1(n154), .A2(n266), .B1(n528), .B2(n97), .ZN(n428) );
  OAI22_X2 U160 ( .A1(n155), .A2(n266), .B1(n528), .B2(n96), .ZN(n429) );
  NAND3_X2 U161 ( .A1(n230), .A2(n229), .A3(n265), .ZN(n266) );
  NAND2_X2 U164 ( .A1(n561), .A2(n499), .ZN(n203) );
  NAND2_X2 U165 ( .A1(n499), .A2(n205), .ZN(n211) );
  NAND2_X2 U166 ( .A1(n559), .A2(n499), .ZN(n229) );
  OAI22_X2 U167 ( .A1(n156), .A2(n267), .B1(n535), .B2(n95), .ZN(n430) );
  NAND3_X2 U168 ( .A1(n251), .A2(n194), .A3(n230), .ZN(n267) );
  OAI22_X2 U169 ( .A1(n544), .A2(n157), .B1(n269), .B2(n94), .ZN(n431) );
  OAI22_X2 U170 ( .A1(n544), .A2(n158), .B1(n269), .B2(n93), .ZN(n432) );
  OAI22_X2 U171 ( .A1(n544), .A2(n159), .B1(n269), .B2(n92), .ZN(n433) );
  OAI22_X2 U173 ( .A1(n543), .A2(n151), .B1(n271), .B2(n91), .ZN(n434) );
  OAI22_X2 U174 ( .A1(n543), .A2(n153), .B1(n271), .B2(n90), .ZN(n435) );
  OAI22_X2 U175 ( .A1(n543), .A2(n154), .B1(n271), .B2(n89), .ZN(n436) );
  NAND4_X2 U177 ( .A1(n272), .A2(n551), .A3(n273), .A4(n164), .ZN(n270) );
  NAND2_X2 U179 ( .A1(WriteBus[75]), .A2(n274), .ZN(n275) );
  NAND2_X2 U181 ( .A1(WriteBus[76]), .A2(n274), .ZN(n276) );
  NAND2_X2 U183 ( .A1(WriteBus[77]), .A2(n274), .ZN(n277) );
  NAND2_X2 U185 ( .A1(WriteBus[78]), .A2(n274), .ZN(n278) );
  NAND2_X2 U187 ( .A1(WriteBus[79]), .A2(n274), .ZN(n279) );
  OAI22_X2 U189 ( .A1(n151), .A2(n282), .B1(n531), .B2(n88), .ZN(n442) );
  NAND3_X2 U190 ( .A1(n169), .A2(n268), .A3(n280), .ZN(n282) );
  OAI22_X2 U191 ( .A1(n153), .A2(n283), .B1(n530), .B2(n87), .ZN(n443) );
  NAND3_X2 U192 ( .A1(n237), .A2(n210), .A3(n169), .ZN(n283) );
  NAND2_X2 U195 ( .A1(WriteBus[82]), .A2(n286), .ZN(n287) );
  NAND2_X2 U197 ( .A1(WriteBus[83]), .A2(n286), .ZN(n288) );
  NAND2_X2 U199 ( .A1(WriteBus[84]), .A2(n286), .ZN(n289) );
  NAND2_X2 U201 ( .A1(WriteBus[85]), .A2(n286), .ZN(n290) );
  NAND2_X2 U203 ( .A1(WriteBus[86]), .A2(n286), .ZN(n291) );
  NAND2_X2 U205 ( .A1(WriteBus[87]), .A2(n286), .ZN(n292) );
  NAND2_X2 U208 ( .A1(n162), .A2(n167), .ZN(n295) );
  NAND3_X2 U209 ( .A1(n263), .A2(n296), .A3(n273), .ZN(n294) );
  NAND2_X2 U211 ( .A1(WriteBus[88]), .A2(n297), .ZN(n298) );
  NAND4_X2 U212 ( .A1(n280), .A2(n284), .A3(n281), .A4(n268), .ZN(n297) );
  NAND2_X2 U213 ( .A1(n571), .A2(n499), .ZN(n268) );
  NAND2_X2 U214 ( .A1(n558), .A2(n499), .ZN(n281) );
  NOR2_X2 U215 ( .A1(n188), .A2(n299), .ZN(n284) );
  NAND2_X2 U217 ( .A1(WriteBus[89]), .A2(n300), .ZN(n301) );
  NAND2_X2 U219 ( .A1(WriteBus[90]), .A2(n300), .ZN(n302) );
  NAND2_X2 U221 ( .A1(WriteBus[91]), .A2(n300), .ZN(n303) );
  NAND2_X2 U223 ( .A1(WriteBus[92]), .A2(n300), .ZN(n304) );
  NAND2_X2 U225 ( .A1(WriteBus[93]), .A2(n300), .ZN(n305) );
  NAND2_X2 U227 ( .A1(WriteBus[94]), .A2(n300), .ZN(n306) );
  NOR4_X2 U229 ( .A1(n308), .A2(n566), .A3(n568), .A4(n262), .ZN(n307) );
  NAND2_X2 U231 ( .A1(WriteBus[95]), .A2(n309), .ZN(n310) );
  NOR3_X2 U233 ( .A1(n568), .A2(n299), .A3(n547), .ZN(n272) );
  NAND2_X2 U235 ( .A1(WriteBus[96]), .A2(n313), .ZN(n314) );
  NAND2_X2 U237 ( .A1(WriteBus[97]), .A2(n313), .ZN(n315) );
  NAND2_X2 U239 ( .A1(WriteBus[98]), .A2(n313), .ZN(n316) );
  NAND2_X2 U241 ( .A1(WriteBus[99]), .A2(n313), .ZN(n317) );
  NAND2_X2 U243 ( .A1(WriteBus[100]), .A2(n313), .ZN(n318) );
  NAND2_X2 U246 ( .A1(WriteBus[101]), .A2(n320), .ZN(n321) );
  NAND4_X2 U247 ( .A1(n246), .A2(n322), .A3(n323), .A4(n251), .ZN(n320) );
  NOR2_X2 U248 ( .A1(n285), .A2(n299), .ZN(n323) );
  NOR2_X2 U249 ( .A1(n273), .A2(n500), .ZN(n285) );
  NAND2_X2 U251 ( .A1(n324), .A2(n189), .ZN(n233) );
  OAI22_X2 U252 ( .A1(n553), .A2(n158), .B1(n325), .B2(n86), .ZN(n464) );
  OAI22_X2 U253 ( .A1(n553), .A2(n159), .B1(n325), .B2(n85), .ZN(n465) );
  OAI22_X2 U255 ( .A1(n552), .A2(n151), .B1(n327), .B2(n84), .ZN(n466) );
  OAI22_X2 U256 ( .A1(n552), .A2(n153), .B1(n327), .B2(n83), .ZN(n467) );
  OAI22_X2 U257 ( .A1(n552), .A2(n154), .B1(n327), .B2(n82), .ZN(n468) );
  OAI22_X2 U258 ( .A1(n552), .A2(n155), .B1(n327), .B2(n81), .ZN(n469) );
  NAND4_X2 U260 ( .A1(n311), .A2(n328), .A3(n273), .A4(n565), .ZN(n326) );
  OAI22_X2 U261 ( .A1(n156), .A2(n329), .B1(n541), .B2(n80), .ZN(n470) );
  NOR3_X2 U263 ( .A1(n569), .A2(n308), .A3(n568), .ZN(n330) );
  OAI22_X2 U264 ( .A1(n157), .A2(n545), .B1(n332), .B2(n79), .ZN(n471) );
  OAI22_X2 U265 ( .A1(n158), .A2(n545), .B1(n332), .B2(n78), .ZN(n472) );
  OAI22_X2 U266 ( .A1(n159), .A2(n545), .B1(n332), .B2(n77), .ZN(n473) );
  NOR2_X2 U267 ( .A1(n333), .A2(n188), .ZN(n332) );
  NAND2_X2 U268 ( .A1(n246), .A2(n546), .ZN(n188) );
  OAI22_X2 U270 ( .A1(n151), .A2(n336), .B1(n542), .B2(n76), .ZN(n474) );
  OAI22_X2 U271 ( .A1(n153), .A2(n336), .B1(n542), .B2(n75), .ZN(n475) );
  OAI22_X2 U272 ( .A1(n154), .A2(n336), .B1(n542), .B2(n74), .ZN(n476) );
  NAND3_X2 U273 ( .A1(n548), .A2(n260), .A3(n337), .ZN(n336) );
  NOR3_X2 U274 ( .A1(n335), .A2(n334), .A3(n299), .ZN(n337) );
  NOR2_X2 U275 ( .A1(n191), .A2(n500), .ZN(n299) );
  NOR2_X2 U276 ( .A1(n331), .A2(n500), .ZN(n334) );
  NOR2_X2 U277 ( .A1(n565), .A2(n500), .ZN(n335) );
  NOR3_X2 U280 ( .A1(n172), .A2(n567), .A3(n560), .ZN(n338) );
  NAND2_X2 U281 ( .A1(n324), .A2(n167), .ZN(n206) );
  NOR2_X2 U282 ( .A1(n180), .A2(n559), .ZN(n324) );
  NAND2_X2 U284 ( .A1(WriteBus[115]), .A2(n340), .ZN(n341) );
  NAND2_X2 U286 ( .A1(WriteBus[116]), .A2(n340), .ZN(n342) );
  NAND2_X2 U288 ( .A1(WriteBus[117]), .A2(n340), .ZN(n343) );
  NAND2_X2 U290 ( .A1(WriteBus[118]), .A2(n340), .ZN(n344) );
  NAND2_X2 U292 ( .A1(WriteBus[119]), .A2(n340), .ZN(n345) );
  NOR2_X2 U294 ( .A1(n247), .A2(n308), .ZN(n346) );
  NOR4_X2 U295 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(n308) );
  NAND2_X2 U297 ( .A1(WriteBus[120]), .A2(n347), .ZN(n348) );
  NOR2_X2 U300 ( .A1(n247), .A2(n569), .ZN(n349) );
  NOR3_X2 U301 ( .A1(n180), .A2(n562), .A3(n181), .ZN(n311) );
  NAND4_X2 U302 ( .A1(n557), .A2(n167), .A3(n350), .A4(n260), .ZN(n181) );
  NOR2_X2 U303 ( .A1(n559), .A2(n558), .ZN(n350) );
  NAND3_X2 U304 ( .A1(n339), .A2(n193), .A3(n162), .ZN(n171) );
  NOR2_X2 U305 ( .A1(n570), .A2(n561), .ZN(n162) );
  NAND2_X2 U306 ( .A1(n190), .A2(n263), .ZN(n180) );
  OAI22_X2 U307 ( .A1(n153), .A2(n352), .B1(n550), .B2(n73), .ZN(n483) );
  OAI22_X2 U309 ( .A1(n154), .A2(n352), .B1(n550), .B2(n72), .ZN(n484) );
  OAI22_X2 U311 ( .A1(n155), .A2(n352), .B1(n550), .B2(n71), .ZN(n485) );
  OAI22_X2 U313 ( .A1(n156), .A2(n352), .B1(n550), .B2(n70), .ZN(n486) );
  OAI22_X2 U315 ( .A1(n157), .A2(n352), .B1(n550), .B2(n69), .ZN(n487) );
  OAI22_X2 U317 ( .A1(n158), .A2(n352), .B1(n550), .B2(n68), .ZN(n488) );
  OAI22_X2 U319 ( .A1(n159), .A2(n352), .B1(n550), .B2(n67), .ZN(n489) );
  NAND3_X2 U320 ( .A1(n353), .A2(n260), .A3(n280), .ZN(n352) );
  AND3_X2 U321 ( .A1(n194), .A2(n184), .A3(n251), .ZN(n280) );
  NAND2_X2 U322 ( .A1(n499), .A2(n354), .ZN(n251) );
  NAND3_X2 U323 ( .A1(n163), .A2(n351), .A3(n555), .ZN(n354) );
  NAND2_X2 U324 ( .A1(n164), .A2(n193), .ZN(n205) );
  NAND3_X2 U325 ( .A1(n65), .A2(n64), .A3(n355), .ZN(n164) );
  NAND2_X2 U326 ( .A1(n356), .A2(n355), .ZN(n351) );
  NAND3_X2 U327 ( .A1(n66), .A2(n63), .A3(n356), .ZN(n339) );
  NAND3_X2 U328 ( .A1(n65), .A2(n63), .A3(n357), .ZN(n234) );
  NAND3_X2 U329 ( .A1(n355), .A2(n65), .A3(\sub_63/A[2] ), .ZN(n224) );
  NAND2_X2 U330 ( .A1(n563), .A2(n499), .ZN(n184) );
  NAND3_X2 U331 ( .A1(n66), .A2(n64), .A3(n358), .ZN(n263) );
  NAND3_X2 U333 ( .A1(\sub_63/A[1] ), .A2(n63), .A3(n357), .ZN(n221) );
  NAND3_X2 U334 ( .A1(\sub_63/A[1] ), .A2(n355), .A3(\sub_63/A[2] ), .ZN(n296)
         );
  NOR2_X2 U335 ( .A1(n66), .A2(\sub_63/A[3] ), .ZN(n355) );
  NAND2_X2 U336 ( .A1(\sub_63/A[4] ), .A2(n499), .ZN(n260) );
  NAND3_X2 U338 ( .A1(n189), .A2(n190), .A3(n328), .ZN(n262) );
  NAND3_X2 U339 ( .A1(\sub_63/A[3] ), .A2(\sub_63/A[1] ), .A3(n357), .ZN(n328)
         );
  NAND3_X2 U340 ( .A1(\sub_63/A[0] ), .A2(n64), .A3(n358), .ZN(n190) );
  NAND3_X2 U341 ( .A1(\sub_63/A[3] ), .A2(n66), .A3(n356), .ZN(n189) );
  NAND3_X2 U342 ( .A1(n191), .A2(n273), .A3(n331), .ZN(n247) );
  NAND2_X2 U343 ( .A1(n357), .A2(n358), .ZN(n331) );
  NOR2_X2 U344 ( .A1(n64), .A2(\sub_63/A[0] ), .ZN(n357) );
  NAND3_X2 U345 ( .A1(\sub_63/A[3] ), .A2(\sub_63/A[0] ), .A3(n356), .ZN(n273)
         );
  NOR2_X2 U346 ( .A1(n65), .A2(\sub_63/A[2] ), .ZN(n356) );
  NAND3_X2 U347 ( .A1(\sub_63/A[2] ), .A2(\sub_63/A[0] ), .A3(n358), .ZN(n191)
         );
  NOR2_X2 U348 ( .A1(n63), .A2(\sub_63/A[1] ), .ZN(n358) );
  NAND2_X2 U350 ( .A1(\sub_63/A[0] ), .A2(n549), .ZN(\U7/Z_0 ) );
  NAND2_X2 U351 ( .A1(n499), .A2(n359), .ZN(n136) );
  NOR2_X2 U352 ( .A1(n500), .A2(n359), .ZN(\U6/Z_0 ) );
  NAND4_X2 U353 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(n193) );
  AND2_X1 U416 ( .A1(n204), .A2(n268), .ZN(n230) );
  AND2_X1 U417 ( .A1(n169), .A2(n281), .ZN(n204) );
  AND2_X1 U418 ( .A1(n284), .A2(n540), .ZN(n169) );
  AND2_X1 U420 ( .A1(n312), .A2(n260), .ZN(n246) );
  OR2_X1 U421 ( .A1(n206), .A2(n558), .ZN(n172) );
  AND2_X1 U422 ( .A1(n167), .A2(n339), .ZN(n163) );
  AND2_X1 U423 ( .A1(n224), .A2(n234), .ZN(n167) );
  OR2_X1 U424 ( .A1(\U5/DATA2_3 ), .A2(n136), .ZN(\U7/Z_3 ) );
  OR2_X1 U425 ( .A1(\U5/DATA2_2 ), .A2(n136), .ZN(\U7/Z_2 ) );
  OR2_X1 U426 ( .A1(\U5/DATA2_1 ), .A2(n136), .ZN(\U7/Z_1 ) );
  OR2_X1 U427 ( .A1(n193), .A2(\sub_63/A[4] ), .ZN(n359) );
  DFFR_X2 \WriteBus_reg[81]  ( .D(n443), .CK(clock), .RN(n504), .Q(
        WriteBus[81]), .QN(n87) );
  DFFR_X2 \WriteBus_reg[80]  ( .D(n442), .CK(clock), .RN(n505), .Q(
        WriteBus[80]), .QN(n88) );
  DFFR_X2 \WriteBus_reg[68]  ( .D(n430), .CK(clock), .RN(n506), .Q(
        WriteBus[68]), .QN(n95) );
  DFFR_X2 \WriteBus_reg[48]  ( .D(n410), .CK(clock), .RN(n507), .Q(
        WriteBus[48]), .QN(n102) );
  DFFR_X2 \WriteBus_reg[9]  ( .D(n371), .CK(clock), .RN(n509), .Q(WriteBus[9]), 
        .QN(n120) );
  DFFR_X2 \WriteBus_reg[8]  ( .D(n370), .CK(clock), .RN(n508), .Q(WriteBus[8]), 
        .QN(n121) );
  DFFR_X2 \WriteBus_reg[127]  ( .D(n489), .CK(clock), .RN(n501), .Q(
        WriteBus[127]), .QN(n67) );
  DFFR_X2 \WriteBus_reg[126]  ( .D(n488), .CK(clock), .RN(n501), .Q(
        WriteBus[126]), .QN(n68) );
  DFFR_X2 \WriteBus_reg[125]  ( .D(n487), .CK(clock), .RN(n501), .Q(
        WriteBus[125]), .QN(n69) );
  DFFR_X2 \WriteBus_reg[124]  ( .D(n486), .CK(clock), .RN(n501), .Q(
        WriteBus[124]), .QN(n70) );
  DFFR_X2 \WriteBus_reg[123]  ( .D(n485), .CK(clock), .RN(n501), .Q(
        WriteBus[123]), .QN(n71) );
  DFFR_X2 \WriteBus_reg[122]  ( .D(n484), .CK(clock), .RN(n501), .Q(
        WriteBus[122]), .QN(n72) );
  DFFR_X2 \WriteBus_reg[121]  ( .D(n483), .CK(clock), .RN(n501), .Q(
        WriteBus[121]), .QN(n73) );
  DFFR_X2 \WriteBus_reg[114]  ( .D(n476), .CK(clock), .RN(n502), .Q(
        WriteBus[114]), .QN(n74) );
  DFFR_X2 \WriteBus_reg[113]  ( .D(n475), .CK(clock), .RN(n502), .Q(
        WriteBus[113]), .QN(n75) );
  DFFR_X2 \WriteBus_reg[112]  ( .D(n474), .CK(clock), .RN(n502), .Q(
        WriteBus[112]), .QN(n76) );
  DFFR_X2 \WriteBus_reg[111]  ( .D(n473), .CK(clock), .RN(n502), .Q(
        WriteBus[111]), .QN(n77) );
  DFFR_X2 \WriteBus_reg[110]  ( .D(n472), .CK(clock), .RN(n502), .Q(
        WriteBus[110]), .QN(n78) );
  DFFR_X2 \WriteBus_reg[109]  ( .D(n471), .CK(clock), .RN(n502), .Q(
        WriteBus[109]), .QN(n79) );
  DFFR_X2 \WriteBus_reg[108]  ( .D(n470), .CK(clock), .RN(n502), .Q(
        WriteBus[108]), .QN(n80) );
  DFFR_X2 \WriteBus_reg[107]  ( .D(n469), .CK(clock), .RN(n502), .Q(
        WriteBus[107]), .QN(n81) );
  DFFR_X2 \WriteBus_reg[106]  ( .D(n468), .CK(clock), .RN(n502), .Q(
        WriteBus[106]), .QN(n82) );
  DFFR_X2 \WriteBus_reg[105]  ( .D(n467), .CK(clock), .RN(n503), .Q(
        WriteBus[105]), .QN(n83) );
  DFFR_X2 \WriteBus_reg[104]  ( .D(n466), .CK(clock), .RN(n503), .Q(
        WriteBus[104]), .QN(n84) );
  DFFR_X2 \WriteBus_reg[103]  ( .D(n465), .CK(clock), .RN(n503), .Q(
        WriteBus[103]), .QN(n85) );
  DFFR_X2 \WriteBus_reg[102]  ( .D(n464), .CK(clock), .RN(n503), .Q(
        WriteBus[102]), .QN(n86) );
  DFFR_X2 \WriteBus_reg[74]  ( .D(n436), .CK(clock), .RN(n505), .Q(
        WriteBus[74]), .QN(n89) );
  DFFR_X2 \WriteBus_reg[73]  ( .D(n435), .CK(clock), .RN(n505), .Q(
        WriteBus[73]), .QN(n90) );
  DFFR_X2 \WriteBus_reg[72]  ( .D(n434), .CK(clock), .RN(n505), .Q(
        WriteBus[72]), .QN(n91) );
  DFFR_X2 \WriteBus_reg[71]  ( .D(n433), .CK(clock), .RN(n505), .Q(
        WriteBus[71]), .QN(n92) );
  DFFR_X2 \WriteBus_reg[70]  ( .D(n432), .CK(clock), .RN(n505), .Q(
        WriteBus[70]), .QN(n93) );
  DFFR_X2 \WriteBus_reg[69]  ( .D(n431), .CK(clock), .RN(n505), .Q(
        WriteBus[69]), .QN(n94) );
  DFFR_X2 \WriteBus_reg[67]  ( .D(n429), .CK(clock), .RN(n506), .Q(
        WriteBus[67]), .QN(n96) );
  DFFR_X2 \WriteBus_reg[66]  ( .D(n428), .CK(clock), .RN(n506), .Q(
        WriteBus[66]), .QN(n97) );
  DFFR_X2 \WriteBus_reg[65]  ( .D(n427), .CK(clock), .RN(n506), .Q(
        WriteBus[65]), .QN(n98) );
  DFFR_X2 \WriteBus_reg[64]  ( .D(n426), .CK(clock), .RN(n506), .Q(
        WriteBus[64]), .QN(n99) );
  DFFR_X2 \WriteBus_reg[63]  ( .D(n425), .CK(clock), .RN(n506), .Q(
        WriteBus[63]), .QN(n100) );
  DFFR_X2 \WriteBus_reg[62]  ( .D(n424), .CK(clock), .RN(n506), .Q(
        WriteBus[62]), .QN(n101) );
  DFFR_X2 \WriteBus_reg[47]  ( .D(n409), .CK(clock), .RN(n507), .Q(
        WriteBus[47]), .QN(n103) );
  DFFR_X2 \WriteBus_reg[46]  ( .D(n408), .CK(clock), .RN(n507), .Q(
        WriteBus[46]), .QN(n104) );
  DFFR_X2 \WriteBus_reg[45]  ( .D(n407), .CK(clock), .RN(n508), .Q(
        WriteBus[45]), .QN(n105) );
  DFFR_X2 \WriteBus_reg[44]  ( .D(n406), .CK(clock), .RN(n508), .Q(
        WriteBus[44]), .QN(n106) );
  DFFR_X2 \WriteBus_reg[43]  ( .D(n405), .CK(clock), .RN(n508), .Q(
        WriteBus[43]), .QN(n107) );
  DFFR_X2 \WriteBus_reg[42]  ( .D(n404), .CK(clock), .RN(n508), .Q(
        WriteBus[42]), .QN(n108) );
  DFFR_X2 \WriteBus_reg[39]  ( .D(n401), .CK(clock), .RN(n508), .Q(
        WriteBus[39]), .QN(n109) );
  DFFR_X2 \WriteBus_reg[38]  ( .D(n400), .CK(clock), .RN(n508), .Q(
        WriteBus[38]), .QN(n110) );
  DFFR_X2 \WriteBus_reg[37]  ( .D(n399), .CK(clock), .RN(n508), .Q(
        WriteBus[37]), .QN(n111) );
  DFFR_X2 \WriteBus_reg[36]  ( .D(n398), .CK(clock), .RN(n508), .Q(
        WriteBus[36]), .QN(n112) );
  DFFR_X2 \WriteBus_reg[35]  ( .D(n397), .CK(clock), .RN(n508), .Q(
        WriteBus[35]), .QN(n113) );
  DFFR_X2 \WriteBus_reg[34]  ( .D(n396), .CK(clock), .RN(n508), .Q(
        WriteBus[34]), .QN(n114) );
  DFFR_X2 \WriteBus_reg[33]  ( .D(n395), .CK(clock), .RN(n509), .Q(
        WriteBus[33]), .QN(n115) );
  DFFR_X2 \WriteBus_reg[32]  ( .D(n394), .CK(clock), .RN(n509), .Q(
        WriteBus[32]), .QN(n116) );
  DFFR_X2 \WriteBus_reg[31]  ( .D(n393), .CK(clock), .RN(n509), .Q(
        WriteBus[31]), .QN(n117) );
  DFFR_X2 \WriteBus_reg[30]  ( .D(n392), .CK(clock), .RN(n509), .Q(
        WriteBus[30]), .QN(n118) );
  DFFR_X2 \WriteBus_reg[29]  ( .D(n391), .CK(clock), .RN(n509), .Q(
        WriteBus[29]), .QN(n119) );
  DFFR_X2 \WriteBus_reg[7]  ( .D(n369), .CK(clock), .RN(n510), .Q(WriteBus[7]), 
        .QN(n122) );
  DFFR_X2 \WriteBus_reg[6]  ( .D(n368), .CK(clock), .RN(n501), .Q(WriteBus[6]), 
        .QN(n123) );
  DFFR_X2 \WriteBus_reg[5]  ( .D(n367), .CK(clock), .RN(n510), .Q(WriteBus[5]), 
        .QN(n124) );
  DFFR_X2 \WriteBus_reg[4]  ( .D(n366), .CK(clock), .RN(n509), .Q(WriteBus[4]), 
        .QN(n125) );
  DFFR_X2 \WriteBus_reg[3]  ( .D(n365), .CK(clock), .RN(n507), .Q(WriteBus[3]), 
        .QN(n126) );
  DFFR_X2 \WriteBus_reg[2]  ( .D(n364), .CK(clock), .RN(n505), .Q(WriteBus[2]), 
        .QN(n127) );
  DFFR_X2 \WriteBus_reg[1]  ( .D(n363), .CK(clock), .RN(n506), .Q(WriteBus[1]), 
        .QN(n128) );
  DFFR_X2 \WriteBus_reg[0]  ( .D(n362), .CK(clock), .RN(n508), .Q(WriteBus[0]), 
        .QN(n129) );
  DFF_X2 \WriteAddress_reg[15]  ( .D(\add_55/A[15] ), .CK(clock), .Q(
        WriteAddress[15]) );
  DFF_X2 \WriteAddress_reg[14]  ( .D(\add_55/A[14] ), .CK(clock), .Q(
        WriteAddress[14]) );
  DFF_X2 \WriteAddress_reg[13]  ( .D(\add_55/A[13] ), .CK(clock), .Q(
        WriteAddress[13]) );
  DFF_X2 \WriteAddress_reg[12]  ( .D(\add_55/A[12] ), .CK(clock), .Q(
        WriteAddress[12]) );
  DFF_X2 \WriteAddress_reg[11]  ( .D(\add_55/A[11] ), .CK(clock), .Q(
        WriteAddress[11]) );
  DFF_X2 \WriteAddress_reg[10]  ( .D(\add_55/A[10] ), .CK(clock), .Q(
        WriteAddress[10]) );
  DFF_X2 \WriteAddress_reg[9]  ( .D(\add_55/A[9] ), .CK(clock), .Q(
        WriteAddress[9]) );
  DFF_X2 \WriteAddress_reg[8]  ( .D(\add_55/A[8] ), .CK(clock), .Q(
        WriteAddress[8]) );
  DFF_X2 \WriteAddress_reg[7]  ( .D(\add_55/A[7] ), .CK(clock), .Q(
        WriteAddress[7]) );
  DFF_X2 \WriteAddress_reg[6]  ( .D(\add_55/A[6] ), .CK(clock), .Q(
        WriteAddress[6]) );
  DFF_X2 \WriteAddress_reg[5]  ( .D(\add_55/A[5] ), .CK(clock), .Q(
        WriteAddress[5]) );
  DFF_X2 \WriteAddress_reg[4]  ( .D(\add_55/A[4] ), .CK(clock), .Q(
        WriteAddress[4]) );
  DFF_X2 \WriteAddress_reg[3]  ( .D(\add_55/A[3] ), .CK(clock), .Q(
        WriteAddress[3]) );
  DFF_X2 \WriteAddress_reg[2]  ( .D(\add_55/A[2] ), .CK(clock), .Q(
        WriteAddress[2]) );
  DFF_X2 \WriteAddress_reg[1]  ( .D(\add_55/A[1] ), .CK(clock), .Q(
        WriteAddress[1]) );
  DFF_X2 \WriteAddress_reg[0]  ( .D(\add_55/A[0] ), .CK(clock), .Q(
        WriteAddress[0]) );
  DFFR_X2 \next_WriteAddress_reg[0]  ( .D(n361), .CK(clock), .RN(n501), .Q(
        \add_55/A[0] ), .QN(n131) );
  DFFR_X2 WriteEnable_reg ( .D(\U6/Z_0 ), .CK(clock), .RN(n501), .Q(
        WriteEnable) );
  DFFR_X2 \next_WriteAddress_reg[2]  ( .D(n515), .CK(clock), .RN(n511), .Q(
        \add_55/A[2] ) );
  DFFR_X2 \next_WriteAddress_reg[1]  ( .D(n514), .CK(clock), .RN(n511), .Q(
        \add_55/A[1] ) );
  DFFR_X2 \WriteBus_reg[55]  ( .D(n417), .CK(clock), .RN(n507), .Q(
        WriteBus[55]) );
  DFFR_X2 \WriteBus_reg[101]  ( .D(n463), .CK(clock), .RN(n503), .Q(
        WriteBus[101]) );
  DFFR_X2 \WriteBus_reg[120]  ( .D(n482), .CK(clock), .RN(n501), .Q(
        WriteBus[120]) );
  DFFR_X2 \WriteBus_reg[95]  ( .D(n457), .CK(clock), .RN(n503), .Q(
        WriteBus[95]) );
  DFFR_X2 \WriteBus_reg[61]  ( .D(n423), .CK(clock), .RN(n506), .Q(
        WriteBus[61]) );
  DFFR_X2 \WriteBus_reg[60]  ( .D(n422), .CK(clock), .RN(n506), .Q(
        WriteBus[60]) );
  DFFR_X2 \WriteBus_reg[59]  ( .D(n421), .CK(clock), .RN(n506), .Q(
        WriteBus[59]) );
  DFFR_X2 \WriteBus_reg[58]  ( .D(n420), .CK(clock), .RN(n506), .Q(
        WriteBus[58]) );
  DFFR_X2 \WriteBus_reg[57]  ( .D(n419), .CK(clock), .RN(n506), .Q(
        WriteBus[57]) );
  DFFR_X2 \WriteBus_reg[56]  ( .D(n418), .CK(clock), .RN(n507), .Q(
        WriteBus[56]) );
  DFFR_X2 \WriteBus_reg[88]  ( .D(n450), .CK(clock), .RN(n504), .Q(
        WriteBus[88]) );
  DFFR_X2 \WriteBus_reg[119]  ( .D(n481), .CK(clock), .RN(n501), .Q(
        WriteBus[119]) );
  DFFR_X2 \WriteBus_reg[118]  ( .D(n480), .CK(clock), .RN(n501), .Q(
        WriteBus[118]) );
  DFFR_X2 \WriteBus_reg[117]  ( .D(n479), .CK(clock), .RN(n502), .Q(
        WriteBus[117]) );
  DFFR_X2 \WriteBus_reg[116]  ( .D(n478), .CK(clock), .RN(n502), .Q(
        WriteBus[116]) );
  DFFR_X2 \WriteBus_reg[115]  ( .D(n477), .CK(clock), .RN(n502), .Q(
        WriteBus[115]) );
  DFFR_X2 \WriteBus_reg[87]  ( .D(n449), .CK(clock), .RN(n504), .Q(
        WriteBus[87]) );
  DFFR_X2 \WriteBus_reg[86]  ( .D(n448), .CK(clock), .RN(n504), .Q(
        WriteBus[86]) );
  DFFR_X2 \WriteBus_reg[85]  ( .D(n447), .CK(clock), .RN(n504), .Q(
        WriteBus[85]) );
  DFFR_X2 \WriteBus_reg[84]  ( .D(n446), .CK(clock), .RN(n504), .Q(
        WriteBus[84]) );
  DFFR_X2 \WriteBus_reg[83]  ( .D(n445), .CK(clock), .RN(n504), .Q(
        WriteBus[83]) );
  DFFR_X2 \WriteBus_reg[82]  ( .D(n444), .CK(clock), .RN(n504), .Q(
        WriteBus[82]) );
  DFFR_X2 \WriteBus_reg[14]  ( .D(n376), .CK(clock), .RN(n510), .Q(
        WriteBus[14]) );
  DFFR_X2 \WriteBus_reg[13]  ( .D(n375), .CK(clock), .RN(n510), .Q(
        WriteBus[13]) );
  DFFR_X2 \WriteBus_reg[12]  ( .D(n374), .CK(clock), .RN(n510), .Q(
        WriteBus[12]) );
  DFFR_X2 \WriteBus_reg[11]  ( .D(n373), .CK(clock), .RN(n510), .Q(
        WriteBus[11]) );
  DFFR_X2 \WriteBus_reg[10]  ( .D(n372), .CK(clock), .RN(n510), .Q(
        WriteBus[10]) );
  DFFR_X2 \WriteBus_reg[15]  ( .D(n377), .CK(clock), .RN(n510), .Q(
        WriteBus[15]) );
  DFFR_X2 \WriteBus_reg[54]  ( .D(n416), .CK(clock), .RN(n507), .Q(
        WriteBus[54]) );
  DFFR_X2 \WriteBus_reg[53]  ( .D(n415), .CK(clock), .RN(n507), .Q(
        WriteBus[53]) );
  DFFR_X2 \WriteBus_reg[52]  ( .D(n414), .CK(clock), .RN(n507), .Q(
        WriteBus[52]) );
  DFFR_X2 \WriteBus_reg[51]  ( .D(n413), .CK(clock), .RN(n507), .Q(
        WriteBus[51]) );
  DFFR_X2 \WriteBus_reg[50]  ( .D(n412), .CK(clock), .RN(n507), .Q(
        WriteBus[50]) );
  DFFR_X2 \WriteBus_reg[49]  ( .D(n411), .CK(clock), .RN(n507), .Q(
        WriteBus[49]) );
  DFFR_X2 \WriteBus_reg[94]  ( .D(n456), .CK(clock), .RN(n503), .Q(
        WriteBus[94]) );
  DFFR_X2 \WriteBus_reg[93]  ( .D(n455), .CK(clock), .RN(n503), .Q(
        WriteBus[93]) );
  DFFR_X2 \WriteBus_reg[92]  ( .D(n454), .CK(clock), .RN(n504), .Q(
        WriteBus[92]) );
  DFFR_X2 \WriteBus_reg[91]  ( .D(n453), .CK(clock), .RN(n504), .Q(
        WriteBus[91]) );
  DFFR_X2 \WriteBus_reg[90]  ( .D(n452), .CK(clock), .RN(n504), .Q(
        WriteBus[90]) );
  DFFR_X2 \WriteBus_reg[89]  ( .D(n451), .CK(clock), .RN(n504), .Q(
        WriteBus[89]) );
  DFFR_X2 \WriteBus_reg[98]  ( .D(n460), .CK(clock), .RN(n503), .Q(
        WriteBus[98]) );
  DFFR_X2 \WriteBus_reg[100]  ( .D(n462), .CK(clock), .RN(n503), .Q(
        WriteBus[100]) );
  DFFR_X2 \WriteBus_reg[99]  ( .D(n461), .CK(clock), .RN(n503), .Q(
        WriteBus[99]) );
  DFFR_X2 \WriteBus_reg[97]  ( .D(n459), .CK(clock), .RN(n507), .Q(
        WriteBus[97]) );
  DFFR_X2 \WriteBus_reg[96]  ( .D(n458), .CK(clock), .RN(n503), .Q(
        WriteBus[96]) );
  DFFR_X2 \WriteBus_reg[23]  ( .D(n385), .CK(clock), .RN(n509), .Q(
        WriteBus[23]) );
  DFFR_X2 \WriteBus_reg[22]  ( .D(n384), .CK(clock), .RN(n509), .Q(
        WriteBus[22]) );
  DFFR_X2 \WriteBus_reg[79]  ( .D(n441), .CK(clock), .RN(n505), .Q(
        WriteBus[79]) );
  DFFR_X2 \WriteBus_reg[78]  ( .D(n440), .CK(clock), .RN(n505), .Q(
        WriteBus[78]) );
  DFFR_X2 \WriteBus_reg[77]  ( .D(n439), .CK(clock), .RN(n505), .Q(
        WriteBus[77]) );
  DFFR_X2 \WriteBus_reg[76]  ( .D(n438), .CK(clock), .RN(n505), .Q(
        WriteBus[76]) );
  DFFR_X2 \WriteBus_reg[75]  ( .D(n437), .CK(clock), .RN(n505), .Q(
        WriteBus[75]) );
  DFFR_X2 \WriteBus_reg[28]  ( .D(n390), .CK(clock), .RN(n509), .Q(
        WriteBus[28]) );
  DFFR_X2 \WriteBus_reg[27]  ( .D(n389), .CK(clock), .RN(n509), .Q(
        WriteBus[27]) );
  DFFR_X2 \WriteBus_reg[26]  ( .D(n388), .CK(clock), .RN(n509), .Q(
        WriteBus[26]) );
  DFFR_X2 \WriteBus_reg[25]  ( .D(n387), .CK(clock), .RN(n509), .Q(
        WriteBus[25]) );
  DFFR_X2 \WriteBus_reg[24]  ( .D(n386), .CK(clock), .RN(n509), .Q(
        WriteBus[24]) );
  DFFR_X2 \WriteBus_reg[21]  ( .D(n383), .CK(clock), .RN(n510), .Q(
        WriteBus[21]) );
  DFFR_X2 \WriteBus_reg[20]  ( .D(n382), .CK(clock), .RN(n510), .Q(
        WriteBus[20]) );
  DFFR_X2 \WriteBus_reg[19]  ( .D(n381), .CK(clock), .RN(n510), .Q(
        WriteBus[19]) );
  DFFR_X2 \WriteBus_reg[18]  ( .D(n380), .CK(clock), .RN(n510), .Q(
        WriteBus[18]) );
  DFFR_X2 \WriteBus_reg[17]  ( .D(n379), .CK(clock), .RN(n510), .Q(
        WriteBus[17]) );
  DFFR_X2 \WriteBus_reg[16]  ( .D(n378), .CK(clock), .RN(n510), .Q(
        WriteBus[16]) );
  DFFR_X2 \WriteBus_reg[41]  ( .D(n403), .CK(clock), .RN(n508), .Q(
        WriteBus[41]) );
  DFFR_X2 \WriteBus_reg[40]  ( .D(n402), .CK(clock), .RN(n508), .Q(
        WriteBus[40]) );
  DFFR_X2 \next_WriteAddress_reg[13]  ( .D(n526), .CK(clock), .RN(n504), .Q(
        \add_55/A[13] ) );
  DFFR_X2 \next_WriteAddress_reg[14]  ( .D(n495), .CK(clock), .RN(n511), .Q(
        \add_55/A[14] ) );
  DFFR_X2 \next_WriteAddress_reg[15]  ( .D(n360), .CK(clock), .RN(n501), .Q(
        \add_55/A[15] ), .QN(n130) );
  OAI22_X1 U4 ( .A1(n136), .A2(n131), .B1(\add_55/A[0] ), .B2(n490), .ZN(n361)
         );
  AND2_X2 U6 ( .A1(\add_55/A[13] ), .A2(n491), .ZN(n492) );
  XOR2_X1 U7 ( .A(\add_55/A[3] ), .B(\add_55/carry[3] ), .Z(\U4/DATA1_3 ) );
  AND2_X2 U8 ( .A1(\add_55/A[3] ), .A2(\add_55/carry[3] ), .ZN(n494) );
  XOR2_X1 U9 ( .A(\add_55/A[9] ), .B(\add_55/carry[9] ), .Z(\U4/DATA1_9 ) );
  AND2_X2 U10 ( .A1(\add_55/A[9] ), .A2(\add_55/carry[9] ), .ZN(n493) );
  INV_X2 U11 ( .A(n135), .ZN(n513) );
  OR2_X4 U12 ( .A1(n500), .A2(n549), .ZN(n490) );
  AND2_X2 U13 ( .A1(\add_55/A[12] ), .A2(\add_55/carry[12] ), .ZN(n491) );
  NAND2_X2 U14 ( .A1(n496), .A2(n497), .ZN(n495) );
  XOR2_X1 U15 ( .A(\add_55/A[13] ), .B(n491), .Z(\U4/DATA1_13 ) );
  XOR2_X1 U16 ( .A(\add_55/A[12] ), .B(\add_55/carry[12] ), .Z(\U4/DATA1_12 )
         );
  NAND2_X2 U17 ( .A1(\U4/DATA1_14 ), .A2(n498), .ZN(n496) );
  NAND2_X2 U18 ( .A1(\add_55/A[14] ), .A2(n549), .ZN(n497) );
  INV_X4 U19 ( .A(n512), .ZN(n506) );
  INV_X4 U20 ( .A(n512), .ZN(n505) );
  INV_X4 U21 ( .A(n512), .ZN(n504) );
  INV_X4 U22 ( .A(n512), .ZN(n507) );
  INV_X4 U38 ( .A(n512), .ZN(n503) );
  INV_X4 U39 ( .A(n512), .ZN(n502) );
  INV_X4 U41 ( .A(n512), .ZN(n511) );
  INV_X4 U43 ( .A(n512), .ZN(n510) );
  INV_X4 U45 ( .A(n512), .ZN(n509) );
  INV_X4 U47 ( .A(n512), .ZN(n508) );
  NAND2_X2 U49 ( .A1(n280), .A2(n204), .ZN(n274) );
  INV_X4 U51 ( .A(n512), .ZN(n501) );
  INV_X4 U54 ( .A(reset_n), .ZN(n512) );
  OAI21_X2 U56 ( .B1(n560), .B2(n206), .A(n499), .ZN(n210) );
  OAI211_X2 U57 ( .C1(n202), .C2(n500), .A(n203), .B(n204), .ZN(n195) );
  OAI211_X2 U59 ( .C1(n218), .C2(n500), .A(n211), .B(n204), .ZN(n212) );
  AOI21_X2 U61 ( .B1(n161), .B2(n556), .A(n500), .ZN(n225) );
  AOI21_X2 U63 ( .B1(n499), .B2(n569), .A(n335), .ZN(n312) );
  INV_X4 U65 ( .A(n500), .ZN(n499) );
  OAI211_X2 U67 ( .C1(n245), .C2(n500), .A(n237), .B(n246), .ZN(n238) );
  OAI211_X2 U69 ( .C1(n179), .C2(n500), .A(n546), .B(n540), .ZN(n173) );
  AOI211_X2 U71 ( .C1(n499), .C2(n570), .A(n554), .B(n187), .ZN(n265) );
  OAI21_X2 U73 ( .B1(n228), .B2(n233), .A(n499), .ZN(n232) );
  OAI21_X2 U76 ( .B1(n568), .B2(n326), .A(n499), .ZN(n327) );
  OAI21_X2 U78 ( .B1(n163), .B2(n500), .A(n203), .ZN(n187) );
  OAI21_X2 U80 ( .B1(n566), .B2(n326), .A(n499), .ZN(n325) );
  AOI21_X2 U82 ( .B1(n312), .B2(n311), .A(n500), .ZN(n319) );
  OAI21_X2 U84 ( .B1(n564), .B2(n205), .A(n499), .ZN(n237) );
  INV_X4 U86 ( .A(n136), .ZN(n549) );
  OAI21_X2 U103 ( .B1(n571), .B2(n270), .A(n499), .ZN(n269) );
  OAI21_X2 U105 ( .B1(n563), .B2(n270), .A(n499), .ZN(n271) );
  OAI21_X2 U107 ( .B1(n559), .B2(n570), .A(n499), .ZN(n194) );
  OAI21_X2 U116 ( .B1(n570), .B2(n233), .A(n499), .ZN(n322) );
  INV_X4 U120 ( .A(n490), .ZN(n498) );
  INV_X4 U121 ( .A(StartIn), .ZN(n500) );
  OAI211_X2 U123 ( .C1(n307), .C2(n500), .A(n260), .B(n280), .ZN(n300) );
  AOI21_X2 U125 ( .B1(n311), .B2(n346), .A(n500), .ZN(n340) );
  NAND4_X2 U127 ( .A1(n284), .A2(n293), .A3(n237), .A4(n268), .ZN(n286) );
  OAI21_X2 U129 ( .B1(n294), .B2(n295), .A(n499), .ZN(n293) );
  OAI21_X2 U131 ( .B1(n247), .B2(n262), .A(n499), .ZN(n353) );
  AOI211_X2 U133 ( .C1(n499), .C2(n186), .A(n187), .B(n188), .ZN(n185) );
  OAI21_X2 U135 ( .B1(n338), .B2(n500), .A(n237), .ZN(n333) );
  OAI211_X2 U138 ( .C1(n259), .C2(n500), .A(n251), .B(n260), .ZN(n252) );
  OAI21_X2 U139 ( .B1(n500), .B2(n193), .A(n194), .ZN(n192) );
  OAI21_X2 U141 ( .B1(n225), .B2(n151), .A(n226), .ZN(n402) );
  OAI21_X2 U143 ( .B1(n225), .B2(n153), .A(n227), .ZN(n403) );
  OAI21_X2 U145 ( .B1(n151), .B2(n195), .A(n196), .ZN(n378) );
  OAI21_X2 U147 ( .B1(n153), .B2(n195), .A(n197), .ZN(n379) );
  OAI21_X2 U149 ( .B1(n154), .B2(n195), .A(n198), .ZN(n380) );
  OAI21_X2 U151 ( .B1(n155), .B2(n195), .A(n199), .ZN(n381) );
  OAI21_X2 U162 ( .B1(n156), .B2(n195), .A(n200), .ZN(n382) );
  OAI21_X2 U163 ( .B1(n157), .B2(n195), .A(n201), .ZN(n383) );
  OAI21_X2 U172 ( .B1(n151), .B2(n212), .A(n213), .ZN(n386) );
  OAI21_X2 U176 ( .B1(n153), .B2(n212), .A(n214), .ZN(n387) );
  OAI21_X2 U178 ( .B1(n154), .B2(n212), .A(n215), .ZN(n388) );
  OAI21_X2 U180 ( .B1(n155), .B2(n212), .A(n216), .ZN(n389) );
  OAI21_X2 U182 ( .B1(n156), .B2(n212), .A(n217), .ZN(n390) );
  OAI21_X2 U184 ( .B1(n513), .B2(n130), .A(n133), .ZN(n360) );
  OAI21_X2 U186 ( .B1(\add_55/carry[15] ), .B2(n500), .A(n136), .ZN(n135) );
  AOI22_X2 U188 ( .A1(\U4/DATA1_13 ), .A2(n498), .B1(\add_55/A[13] ), .B2(n549), .ZN(n138) );
  AOI22_X2 U193 ( .A1(\U4/DATA1_12 ), .A2(n498), .B1(\add_55/A[12] ), .B2(n549), .ZN(n139) );
  AOI22_X2 U194 ( .A1(\U4/DATA1_11 ), .A2(n498), .B1(\add_55/A[11] ), .B2(n549), .ZN(n140) );
  AOI22_X2 U196 ( .A1(\U4/DATA1_10 ), .A2(n498), .B1(\add_55/A[10] ), .B2(n549), .ZN(n141) );
  AOI22_X2 U198 ( .A1(\U4/DATA1_9 ), .A2(n498), .B1(\add_55/A[9] ), .B2(n549), 
        .ZN(n142) );
  OAI21_X2 U200 ( .B1(n171), .B2(n172), .A(n499), .ZN(n170) );
  OAI21_X2 U202 ( .B1(n561), .B2(n172), .A(n499), .ZN(n236) );
  OAI21_X2 U204 ( .B1(n159), .B2(n182), .A(n183), .ZN(n377) );
  OAI21_X2 U206 ( .B1(n347), .B2(n151), .A(n348), .ZN(n482) );
  AOI21_X2 U207 ( .B1(n311), .B2(n349), .A(n500), .ZN(n347) );
  OAI211_X2 U210 ( .C1(n330), .C2(n500), .A(n260), .B(n548), .ZN(n329) );
  OAI21_X2 U216 ( .B1(n154), .B2(n173), .A(n174), .ZN(n372) );
  OAI21_X2 U218 ( .B1(n155), .B2(n173), .A(n175), .ZN(n373) );
  OAI21_X2 U220 ( .B1(n156), .B2(n173), .A(n176), .ZN(n374) );
  OAI21_X2 U222 ( .B1(n157), .B2(n173), .A(n177), .ZN(n375) );
  OAI21_X2 U224 ( .B1(n158), .B2(n173), .A(n178), .ZN(n376) );
  OAI21_X2 U226 ( .B1(n158), .B2(n207), .A(n208), .ZN(n384) );
  OAI21_X2 U228 ( .B1(n159), .B2(n207), .A(n209), .ZN(n385) );
  OAI21_X2 U230 ( .B1(n153), .B2(n238), .A(n239), .ZN(n411) );
  OAI21_X2 U232 ( .B1(n154), .B2(n238), .A(n240), .ZN(n412) );
  OAI21_X2 U234 ( .B1(n155), .B2(n238), .A(n241), .ZN(n413) );
  OAI21_X2 U236 ( .B1(n156), .B2(n238), .A(n242), .ZN(n414) );
  OAI21_X2 U238 ( .B1(n157), .B2(n238), .A(n243), .ZN(n415) );
  OAI21_X2 U240 ( .B1(n158), .B2(n238), .A(n244), .ZN(n416) );
  OAI21_X2 U242 ( .B1(n155), .B2(n274), .A(n275), .ZN(n437) );
  OAI21_X2 U244 ( .B1(n156), .B2(n274), .A(n276), .ZN(n438) );
  OAI21_X2 U245 ( .B1(n157), .B2(n274), .A(n277), .ZN(n439) );
  OAI21_X2 U250 ( .B1(n158), .B2(n274), .A(n278), .ZN(n440) );
  OAI21_X2 U254 ( .B1(n159), .B2(n274), .A(n279), .ZN(n441) );
  OAI21_X2 U259 ( .B1(n154), .B2(n286), .A(n287), .ZN(n444) );
  OAI21_X2 U262 ( .B1(n155), .B2(n286), .A(n288), .ZN(n445) );
  OAI21_X2 U269 ( .B1(n156), .B2(n286), .A(n289), .ZN(n446) );
  OAI21_X2 U278 ( .B1(n157), .B2(n286), .A(n290), .ZN(n447) );
  OAI21_X2 U279 ( .B1(n158), .B2(n286), .A(n291), .ZN(n448) );
  OAI21_X2 U283 ( .B1(n159), .B2(n286), .A(n292), .ZN(n449) );
  OAI21_X2 U285 ( .B1(n151), .B2(n297), .A(n298), .ZN(n450) );
  OAI21_X2 U287 ( .B1(n153), .B2(n300), .A(n301), .ZN(n451) );
  OAI21_X2 U289 ( .B1(n154), .B2(n300), .A(n302), .ZN(n452) );
  OAI21_X2 U291 ( .B1(n155), .B2(n300), .A(n303), .ZN(n453) );
  OAI21_X2 U293 ( .B1(n156), .B2(n300), .A(n304), .ZN(n454) );
  OAI21_X2 U296 ( .B1(n157), .B2(n300), .A(n305), .ZN(n455) );
  OAI21_X2 U298 ( .B1(n158), .B2(n300), .A(n306), .ZN(n456) );
  OAI21_X2 U299 ( .B1(n309), .B2(n159), .A(n310), .ZN(n457) );
  AOI21_X2 U308 ( .B1(n272), .B2(n311), .A(n500), .ZN(n309) );
  OAI21_X2 U310 ( .B1(n151), .B2(n313), .A(n314), .ZN(n458) );
  OAI21_X2 U312 ( .B1(n153), .B2(n313), .A(n315), .ZN(n459) );
  OAI21_X2 U314 ( .B1(n154), .B2(n313), .A(n316), .ZN(n460) );
  OAI21_X2 U316 ( .B1(n155), .B2(n313), .A(n317), .ZN(n461) );
  OAI21_X2 U318 ( .B1(n156), .B2(n313), .A(n318), .ZN(n462) );
  OAI21_X2 U332 ( .B1(n340), .B2(n155), .A(n341), .ZN(n477) );
  OAI21_X2 U337 ( .B1(n340), .B2(n156), .A(n342), .ZN(n478) );
  OAI21_X2 U349 ( .B1(n340), .B2(n157), .A(n343), .ZN(n479) );
  OAI21_X2 U354 ( .B1(n340), .B2(n158), .A(n344), .ZN(n480) );
  OAI21_X2 U355 ( .B1(n340), .B2(n159), .A(n345), .ZN(n481) );
  AOI22_X2 U356 ( .A1(\U4/DATA1_8 ), .A2(n498), .B1(\add_55/A[8] ), .B2(n549), 
        .ZN(n143) );
  AOI22_X2 U357 ( .A1(\U4/DATA1_7 ), .A2(n498), .B1(\add_55/A[7] ), .B2(n549), 
        .ZN(n144) );
  AOI22_X2 U358 ( .A1(\U4/DATA1_6 ), .A2(n498), .B1(\add_55/A[6] ), .B2(n549), 
        .ZN(n145) );
  AOI22_X2 U359 ( .A1(\U4/DATA1_3 ), .A2(n498), .B1(\add_55/A[3] ), .B2(n549), 
        .ZN(n148) );
  AOI22_X2 U360 ( .A1(\U4/DATA1_2 ), .A2(n498), .B1(\add_55/A[2] ), .B2(n549), 
        .ZN(n149) );
  AOI22_X2 U361 ( .A1(\U4/DATA1_1 ), .A2(n498), .B1(\add_55/A[1] ), .B2(n549), 
        .ZN(n150) );
  NAND2_X2 U362 ( .A1(\U8/DATA1_0 ), .A2(n499), .ZN(n151) );
  NAND2_X2 U363 ( .A1(\U8/DATA1_1 ), .A2(n499), .ZN(n153) );
  NAND2_X2 U364 ( .A1(\U8/DATA1_2 ), .A2(n499), .ZN(n154) );
  NAND2_X2 U365 ( .A1(\U8/DATA1_4 ), .A2(n499), .ZN(n156) );
  NAND2_X2 U366 ( .A1(\U8/DATA1_6 ), .A2(n499), .ZN(n158) );
  NAND2_X2 U367 ( .A1(\U8/DATA1_7 ), .A2(n499), .ZN(n159) );
  OAI21_X2 U368 ( .B1(n159), .B2(n248), .A(n249), .ZN(n417) );
  OAI21_X2 U369 ( .B1(n233), .B2(n247), .A(n499), .ZN(n250) );
  OAI21_X2 U370 ( .B1(n151), .B2(n252), .A(n253), .ZN(n418) );
  OAI21_X2 U371 ( .B1(n153), .B2(n252), .A(n254), .ZN(n419) );
  OAI21_X2 U372 ( .B1(n154), .B2(n252), .A(n255), .ZN(n420) );
  OAI21_X2 U373 ( .B1(n155), .B2(n252), .A(n256), .ZN(n421) );
  OAI21_X2 U374 ( .B1(n156), .B2(n252), .A(n257), .ZN(n422) );
  OAI21_X2 U375 ( .B1(n157), .B2(n252), .A(n258), .ZN(n423) );
  OAI21_X2 U376 ( .B1(n157), .B2(n320), .A(n321), .ZN(n463) );
  NAND2_X2 U377 ( .A1(\U8/DATA1_3 ), .A2(n499), .ZN(n155) );
  NAND2_X2 U378 ( .A1(\U8/DATA1_5 ), .A2(n499), .ZN(n157) );
  AOI22_X2 U379 ( .A1(\U4/DATA1_5 ), .A2(n498), .B1(\add_55/A[5] ), .B2(n549), 
        .ZN(n146) );
  AOI22_X2 U380 ( .A1(\U4/DATA1_4 ), .A2(n498), .B1(\add_55/A[4] ), .B2(n549), 
        .ZN(n147) );
  OR3_X4 U381 ( .A1(n299), .A2(n285), .A3(n319), .ZN(n313) );
  INV_X4 U382 ( .A(n150), .ZN(n514) );
  INV_X4 U383 ( .A(n149), .ZN(n515) );
  INV_X4 U384 ( .A(n148), .ZN(n516) );
  INV_X4 U385 ( .A(n147), .ZN(n517) );
  INV_X4 U386 ( .A(n146), .ZN(n518) );
  INV_X4 U387 ( .A(n145), .ZN(n519) );
  INV_X4 U388 ( .A(n144), .ZN(n520) );
  INV_X4 U389 ( .A(n143), .ZN(n521) );
  INV_X4 U390 ( .A(n142), .ZN(n522) );
  INV_X4 U391 ( .A(n141), .ZN(n523) );
  INV_X4 U392 ( .A(n140), .ZN(n524) );
  INV_X4 U393 ( .A(n139), .ZN(n525) );
  INV_X4 U394 ( .A(n138), .ZN(n526) );
  INV_X4 U395 ( .A(n192), .ZN(n527) );
  INV_X4 U396 ( .A(n266), .ZN(n528) );
  INV_X4 U397 ( .A(n264), .ZN(n529) );
  INV_X4 U398 ( .A(n283), .ZN(n530) );
  INV_X4 U399 ( .A(n282), .ZN(n531) );
  INV_X4 U400 ( .A(n235), .ZN(n532) );
  INV_X4 U401 ( .A(n231), .ZN(n533) );
  INV_X4 U402 ( .A(n168), .ZN(n534) );
  INV_X4 U403 ( .A(n267), .ZN(n535) );
  INV_X4 U404 ( .A(n222), .ZN(n536) );
  INV_X4 U405 ( .A(n219), .ZN(n537) );
  INV_X4 U406 ( .A(n165), .ZN(n538) );
  INV_X4 U407 ( .A(n152), .ZN(n539) );
  INV_X4 U408 ( .A(n285), .ZN(n540) );
  INV_X4 U409 ( .A(n329), .ZN(n541) );
  INV_X4 U410 ( .A(n336), .ZN(n542) );
  INV_X4 U411 ( .A(n271), .ZN(n543) );
  INV_X4 U412 ( .A(n269), .ZN(n544) );
  INV_X4 U413 ( .A(n332), .ZN(n545) );
  INV_X4 U414 ( .A(n334), .ZN(n546) );
  INV_X4 U415 ( .A(n312), .ZN(n547) );
  INV_X4 U419 ( .A(n333), .ZN(n548) );
  INV_X4 U428 ( .A(n352), .ZN(n550) );
  INV_X4 U429 ( .A(n181), .ZN(n551) );
  INV_X4 U430 ( .A(n327), .ZN(n552) );
  INV_X4 U431 ( .A(n325), .ZN(n553) );
  INV_X4 U432 ( .A(n211), .ZN(n554) );
  INV_X4 U433 ( .A(n205), .ZN(n555) );
  INV_X4 U434 ( .A(n228), .ZN(n556) );
  INV_X4 U435 ( .A(n171), .ZN(n557) );
  INV_X4 U436 ( .A(n189), .ZN(n558) );
  INV_X4 U437 ( .A(n296), .ZN(n559) );
  INV_X4 U438 ( .A(n162), .ZN(n560) );
  INV_X4 U439 ( .A(n351), .ZN(n561) );
  INV_X4 U440 ( .A(n164), .ZN(n562) );
  INV_X4 U441 ( .A(n263), .ZN(n563) );
  INV_X4 U442 ( .A(n339), .ZN(n564) );
  INV_X4 U443 ( .A(n308), .ZN(n565) );
  INV_X4 U444 ( .A(n191), .ZN(n566) );
  INV_X4 U445 ( .A(n273), .ZN(n567) );
  INV_X4 U446 ( .A(n331), .ZN(n568) );
  INV_X4 U447 ( .A(n328), .ZN(n569) );
  INV_X4 U448 ( .A(n221), .ZN(n570) );
  INV_X4 U449 ( .A(n190), .ZN(n571) );
endmodule


module Output_top ( clock, reset_n, start, CdfMin, divisor, M2SP_ReadBus, 
        M2SP_ReadAddress, M3SP_ReadBus, M3SP_ReadAddress, WriteEnable, 
        Output_MEMBus, Output_MEMAddress, done, output_base_offset );
  input [19:0] CdfMin;
  input [19:0] divisor;
  input [19:0] M2SP_ReadBus;
  output [15:0] M2SP_ReadAddress;
  input [127:0] M3SP_ReadBus;
  output [15:0] M3SP_ReadAddress;
  output [127:0] Output_MEMBus;
  output [15:0] Output_MEMAddress;
  input clock, reset_n, start, output_base_offset;
  output WriteEnable, done;
  wire   start_to_stage_two, start_to_stage_three, start_to_stage_four,
         start_to_stage_five, n15, n16;
  wire   [19:0] DataToStageThree;
  wire   [27:0] DataToStageFour;
  wire   [7:0] result;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  Output_Fetch_MEM stage1 ( .clock(clock), .reset_n(n15), .start(start), 
        .ReadBus(M3SP_ReadBus), .ReadAddress(M3SP_ReadAddress), .DataOut({
        M2SP_ReadAddress[15], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, M2SP_ReadAddress[7:0]}), .StartOut(
        start_to_stage_two), .output_base_offset(output_base_offset), .done(
        done) );
  Output_Fetch_Cdf stage2 ( .clock(clock), .reset_n(n15), .ReadBus(
        M2SP_ReadBus), .DataOut(DataToStageThree), .StartIn(start_to_stage_two), .StartOut(start_to_stage_three) );
  Output_TopExpression stage3 ( .clock(clock), .reset_n(n15), .DataIn(
        DataToStageThree), .CdfMin(CdfMin), .StartIn(start_to_stage_three), 
        .StartOut(start_to_stage_four), .DataOut(DataToStageFour) );
  Output_Result stage4 ( .clock(clock), .reset_n(n15), .DataIn(DataToStageFour), .StartIn(start_to_stage_four), .Divisor(divisor), .StartOut(
        start_to_stage_five), .DataOut(result) );
  Output_Store stage5 ( .clock(clock), .reset_n(n15), .StartIn(
        start_to_stage_five), .ResultIn(result), .WriteBus(Output_MEMBus), 
        .WriteAddress(Output_MEMAddress), .WriteEnable(WriteEnable), 
        .output_base_offset(output_base_offset) );
  INV_X4 U1 ( .A(1'b1), .ZN(M2SP_ReadAddress[8]) );
  INV_X4 U3 ( .A(1'b1), .ZN(M2SP_ReadAddress[9]) );
  INV_X4 U5 ( .A(1'b1), .ZN(M2SP_ReadAddress[10]) );
  INV_X4 U7 ( .A(1'b1), .ZN(M2SP_ReadAddress[11]) );
  INV_X4 U9 ( .A(1'b1), .ZN(M2SP_ReadAddress[12]) );
  INV_X4 U11 ( .A(1'b1), .ZN(M2SP_ReadAddress[13]) );
  INV_X4 U13 ( .A(1'b1), .ZN(M2SP_ReadAddress[14]) );
  INV_X4 U15 ( .A(n16), .ZN(n15) );
  INV_X4 U16 ( .A(reset_n), .ZN(n16) );
endmodule


module Controllor ( clock, reset_n, start, output_start, input_start, 
        input_done, output_done, Cdf_Min, Cdf_Min_Out, Divisor, 
        output_base_offset, input_base_offset, cdf_valid );
  input [19:0] Cdf_Min;
  output [19:0] Cdf_Min_Out;
  output [19:0] Divisor;
  input clock, reset_n, start, input_done, output_done, cdf_valid;
  output output_start, input_start, output_base_offset, input_base_offset;
  wire   \U3/U1/Z_0 , \U15/Z_1 , \U15/Z_2 , \U15/Z_3 , \U15/Z_4 , \U15/Z_5 ,
         \U15/Z_6 , \U15/Z_7 , \U15/Z_8 , \U15/Z_9 , \U15/Z_10 , \U15/Z_11 ,
         \U15/Z_12 , \U15/Z_13 , \U15/Z_14 , \U15/Z_15 , \U15/Z_16 ,
         \U15/Z_17 , \U15/Z_18 , \U15/Z_19 , \U14/DATA1_0 , \U11/DATA1_0 ,
         \U10/DATA2_0 , \r312/DIFF[1] , \r312/DIFF[2] , \r312/DIFF[3] ,
         \r312/DIFF[4] , \r312/DIFF[5] , \r312/DIFF[6] , \r312/DIFF[7] ,
         \r312/DIFF[8] , \r312/DIFF[9] , \r312/DIFF[10] , \r312/DIFF[11] ,
         \r312/DIFF[12] , \r312/DIFF[13] , \r312/DIFF[14] , \r312/DIFF[15] ,
         \r312/DIFF[16] , \r312/DIFF[17] , \r312/DIFF[18] , \r312/DIFF[19] ,
         n24, n25, n26, n27, n30, n31, n33, n34, n37, n39, n41, n42, n43, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n127, n128, n129, n130, n131, n132, n133,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279;
  assign Cdf_Min_Out[0] = \U3/U1/Z_0 ;
  assign Cdf_Min_Out[1] = \U15/Z_1 ;
  assign Cdf_Min_Out[2] = \U15/Z_2 ;
  assign Cdf_Min_Out[3] = \U15/Z_3 ;
  assign Cdf_Min_Out[4] = \U15/Z_4 ;
  assign Cdf_Min_Out[5] = \U15/Z_5 ;
  assign Cdf_Min_Out[6] = \U15/Z_6 ;
  assign Cdf_Min_Out[7] = \U15/Z_7 ;
  assign Cdf_Min_Out[8] = \U15/Z_8 ;
  assign Cdf_Min_Out[9] = \U15/Z_9 ;
  assign Cdf_Min_Out[10] = \U15/Z_10 ;
  assign Cdf_Min_Out[11] = \U15/Z_11 ;
  assign Cdf_Min_Out[12] = \U15/Z_12 ;
  assign Cdf_Min_Out[13] = \U15/Z_13 ;
  assign Cdf_Min_Out[14] = \U15/Z_14 ;
  assign Cdf_Min_Out[15] = \U15/Z_15 ;
  assign Cdf_Min_Out[16] = \U15/Z_16 ;
  assign Cdf_Min_Out[17] = \U15/Z_17 ;
  assign Cdf_Min_Out[18] = \U15/Z_18 ;
  assign Cdf_Min_Out[19] = \U15/Z_19 ;
  assign \U14/DATA1_0  = output_done;
  assign \U11/DATA1_0  = start;
  assign \U10/DATA2_0  = input_done;
  assign Divisor[1] = \r312/DIFF[1] ;
  assign Divisor[2] = \r312/DIFF[2] ;
  assign Divisor[3] = \r312/DIFF[3] ;
  assign Divisor[4] = \r312/DIFF[4] ;
  assign Divisor[5] = \r312/DIFF[5] ;
  assign Divisor[6] = \r312/DIFF[6] ;
  assign Divisor[7] = \r312/DIFF[7] ;
  assign Divisor[8] = \r312/DIFF[8] ;
  assign Divisor[9] = \r312/DIFF[9] ;
  assign Divisor[10] = \r312/DIFF[10] ;
  assign Divisor[11] = \r312/DIFF[11] ;
  assign Divisor[12] = \r312/DIFF[12] ;
  assign Divisor[13] = \r312/DIFF[13] ;
  assign Divisor[14] = \r312/DIFF[14] ;
  assign Divisor[15] = \r312/DIFF[15] ;
  assign Divisor[16] = \r312/DIFF[16] ;
  assign Divisor[17] = \r312/DIFF[17] ;
  assign Divisor[18] = \r312/DIFF[18] ;
  assign Divisor[19] = \r312/DIFF[19] ;

  DFF_X1 RepeatState_reg ( .D(n131), .CK(clock), .QN(n125) );
  DFFR_X1 output_start_reg ( .D(n129), .CK(clock), .RN(reset_n), .Q(
        output_start), .QN(n43) );
  DFFR_X1 input_start_reg ( .D(n130), .CK(clock), .RN(reset_n), .Q(input_start) );
  DFFR_X1 input_base_offset_reg ( .D(n127), .CK(clock), .RN(reset_n), .Q(
        input_base_offset), .QN(n177) );
  DFF_X1 \cdf_min1_reg[0]  ( .D(n123), .CK(cdf_valid), .Q(n217) );
  DFF_X1 \cdf_min1_reg[1]  ( .D(n122), .CK(cdf_valid), .Q(n216) );
  DFF_X1 \cdf_min1_reg[2]  ( .D(n121), .CK(cdf_valid), .Q(n214) );
  DFF_X1 \cdf_min1_reg[3]  ( .D(n120), .CK(cdf_valid), .Q(n215) );
  DFF_X1 \cdf_min1_reg[4]  ( .D(n119), .CK(cdf_valid), .Q(n202) );
  DFF_X1 \cdf_min1_reg[5]  ( .D(n118), .CK(n224), .Q(n203) );
  DFF_X1 \cdf_min1_reg[6]  ( .D(n117), .CK(cdf_valid), .Q(n204) );
  DFF_X1 \cdf_min1_reg[7]  ( .D(n116), .CK(n224), .Q(n205) );
  DFF_X1 \cdf_min1_reg[8]  ( .D(n115), .CK(n224), .Q(n206) );
  DFF_X1 \cdf_min1_reg[9]  ( .D(n114), .CK(cdf_valid), .Q(n207) );
  DFF_X1 \cdf_min1_reg[10]  ( .D(n113), .CK(cdf_valid), .Q(n208) );
  DFF_X1 \cdf_min1_reg[11]  ( .D(n112), .CK(cdf_valid), .Q(n209) );
  DFF_X1 \cdf_min1_reg[12]  ( .D(n111), .CK(cdf_valid), .Q(n210) );
  DFF_X1 \cdf_min1_reg[13]  ( .D(n110), .CK(cdf_valid), .Q(n211) );
  DFF_X1 \cdf_min1_reg[14]  ( .D(n109), .CK(cdf_valid), .Q(n212) );
  DFF_X1 \cdf_min1_reg[15]  ( .D(n108), .CK(cdf_valid), .Q(n213) );
  DFF_X1 \cdf_min1_reg[16]  ( .D(n107), .CK(n224), .Q(n197) );
  DFF_X1 \cdf_min1_reg[17]  ( .D(n106), .CK(n224), .Q(n198) );
  DFF_X1 \cdf_min1_reg[18]  ( .D(n105), .CK(n224), .Q(n199) );
  DFF_X1 \cdf_min1_reg[19]  ( .D(n104), .CK(n224), .Q(n200) );
  DFF_X1 \cdf_min0_reg[19]  ( .D(n103), .CK(cdf_valid), .Q(n181) );
  DFF_X1 \cdf_min0_reg[18]  ( .D(n102), .CK(cdf_valid), .Q(n180) );
  DFF_X1 \cdf_min0_reg[17]  ( .D(n101), .CK(cdf_valid), .Q(n179) );
  DFF_X1 \cdf_min0_reg[16]  ( .D(n100), .CK(cdf_valid), .Q(n178) );
  DFF_X1 \cdf_min0_reg[15]  ( .D(n99), .CK(n224), .Q(n195) );
  DFF_X1 \cdf_min0_reg[14]  ( .D(n98), .CK(cdf_valid), .Q(n194) );
  DFF_X1 \cdf_min0_reg[13]  ( .D(n97), .CK(n224), .Q(n193) );
  DFF_X1 \cdf_min0_reg[12]  ( .D(n96), .CK(cdf_valid), .Q(n192) );
  DFF_X1 \cdf_min0_reg[11]  ( .D(n95), .CK(n224), .Q(n191) );
  DFF_X1 \cdf_min0_reg[10]  ( .D(n94), .CK(n224), .Q(n190) );
  DFF_X1 \cdf_min0_reg[9]  ( .D(n93), .CK(n224), .Q(n189) );
  DFF_X1 \cdf_min0_reg[8]  ( .D(n92), .CK(n224), .Q(n188) );
  DFF_X1 \cdf_min0_reg[7]  ( .D(n91), .CK(n224), .Q(n187) );
  DFF_X1 \cdf_min0_reg[6]  ( .D(n90), .CK(n224), .Q(n186) );
  DFF_X1 \cdf_min0_reg[5]  ( .D(n89), .CK(n224), .Q(n185) );
  DFF_X1 \cdf_min0_reg[4]  ( .D(n88), .CK(n224), .Q(n184) );
  DFF_X1 \cdf_min0_reg[3]  ( .D(n87), .CK(n224), .Q(n183) );
  DFF_X1 \cdf_min0_reg[2]  ( .D(n86), .CK(n224), .Q(n182) );
  DFF_X1 \cdf_min0_reg[1]  ( .D(n85), .CK(n224), .Q(n201) );
  DFF_X1 \cdf_min0_reg[0]  ( .D(n84), .CK(n224), .Q(n196) );
  OR3_X1 U82 ( .A1(n26), .A2(n27), .A3(n37), .ZN(n132) );
  OAI22_X2 U65 ( .A1(n223), .A2(n275), .B1(n24), .B2(n25), .ZN(n127) );
  OAI22_X2 U71 ( .A1(n278), .A2(n43), .B1(\U14/DATA1_0 ), .B2(n31), .ZN(n129)
         );
  NAND3_X2 U72 ( .A1(n31), .A2(n33), .A3(n34), .ZN(n130) );
  NAND2_X2 U74 ( .A1(n274), .A2(n39), .ZN(n131) );
  NAND3_X2 U75 ( .A1(\U14/DATA1_0 ), .A2(n279), .A3(reset_n), .ZN(n39) );
  NAND2_X2 U77 ( .A1(n125), .A2(n26), .ZN(n31) );
  AND3_X2 U83 ( .A1(\U10/DATA2_0 ), .A2(n277), .A3(n42), .ZN(n27) );
  NAND2_X2 U85 ( .A1(n124), .A2(n33), .ZN(n133) );
  NAND3_X2 U86 ( .A1(n124), .A2(n278), .A3(\U11/DATA1_0 ), .ZN(n33) );
  NOR2_X2 U88 ( .A1(n42), .A2(n26), .ZN(n37) );
  NOR2_X2 U89 ( .A1(n42), .A2(n124), .ZN(n26) );
  DFFR_X2 output_base_offset_reg ( .D(n128), .CK(clock), .RN(reset_n), .Q(n176), .QN(n228) );
  DFFR_X2 \State_reg[0]  ( .D(n133), .CK(clock), .RN(reset_n), .Q(n277), .QN(
        n124) );
  DFFR_X2 \State_reg[1]  ( .D(n132), .CK(clock), .RN(reset_n), .QN(n42) );
  BUF_X4 U3 ( .A(n226), .Z(output_base_offset) );
  INV_X1 U4 ( .A(n228), .ZN(n226) );
  INV_X4 U5 ( .A(\U15/Z_2 ), .ZN(n233) );
  INV_X4 U6 ( .A(n234), .ZN(\U15/Z_1 ) );
  NAND2_X2 U7 ( .A1(\U15/Z_12 ), .A2(n255), .ZN(n262) );
  BUF_X4 U8 ( .A(\U3/U1/Z_0 ), .Z(Divisor[0]) );
  NOR2_X1 U9 ( .A1(\U15/Z_7 ), .A2(n244), .ZN(n245) );
  INV_X1 U10 ( .A(\U15/Z_7 ), .ZN(n246) );
  NAND2_X2 U11 ( .A1(n219), .A2(n256), .ZN(n255) );
  OR2_X4 U12 ( .A1(n227), .A2(n201), .ZN(n220) );
  XOR2_X1 U13 ( .A(n233), .B(n231), .Z(\r312/DIFF[2] ) );
  INV_X4 U14 ( .A(n240), .ZN(n218) );
  INV_X4 U15 ( .A(n254), .ZN(n219) );
  INV_X1 U16 ( .A(n254), .ZN(n258) );
  XOR2_X1 U17 ( .A(n237), .B(n239), .Z(\r312/DIFF[3] ) );
  XOR2_X1 U18 ( .A(n238), .B(n236), .Z(\r312/DIFF[4] ) );
  XOR2_X1 U19 ( .A(n246), .B(n248), .Z(\r312/DIFF[7] ) );
  NAND2_X1 U20 ( .A1(n265), .A2(n263), .ZN(\r312/DIFF[13] ) );
  INV_X2 U21 ( .A(\U15/Z_4 ), .ZN(n238) );
  NOR2_X1 U22 ( .A1(\U15/Z_1 ), .A2(\U3/U1/Z_0 ), .ZN(n231) );
  XOR2_X1 U23 ( .A(\U15/Z_1 ), .B(\U3/U1/Z_0 ), .Z(\r312/DIFF[1] ) );
  NAND3_X1 U24 ( .A1(n234), .A2(n233), .A3(n232), .ZN(n235) );
  NAND2_X1 U25 ( .A1(n262), .A2(n259), .ZN(\r312/DIFF[12] ) );
  NAND2_X1 U26 ( .A1(n262), .A2(n261), .ZN(n263) );
  NAND2_X4 U27 ( .A1(n260), .A2(\U15/Z_13 ), .ZN(n265) );
  NOR2_X1 U28 ( .A1(\U15/Z_9 ), .A2(n249), .ZN(n250) );
  OR2_X4 U29 ( .A1(n216), .A2(n228), .ZN(n221) );
  NOR2_X1 U30 ( .A1(\U15/Z_5 ), .A2(n240), .ZN(n241) );
  INV_X1 U31 ( .A(\U15/Z_5 ), .ZN(n242) );
  NOR2_X1 U32 ( .A1(output_base_offset), .A2(n229), .ZN(n230) );
  NOR2_X1 U33 ( .A1(\U15/Z_3 ), .A2(n235), .ZN(n236) );
  NAND2_X2 U34 ( .A1(n220), .A2(n221), .ZN(n234) );
  INV_X1 U35 ( .A(\U15/Z_6 ), .ZN(n243) );
  MUX2_X1 U36 ( .A(n176), .B(n230), .S(n275), .Z(n128) );
  XNOR2_X1 U37 ( .A(n272), .B(\U15/Z_18 ), .ZN(\r312/DIFF[18] ) );
  XNOR2_X2 U38 ( .A(n273), .B(\U15/Z_19 ), .ZN(\r312/DIFF[19] ) );
  OAI21_X1 U39 ( .B1(\U15/Z_15 ), .B2(n266), .A(n268), .ZN(\r312/DIFF[15] ) );
  AOI21_X2 U40 ( .B1(n177), .B2(n26), .A(n27), .ZN(n24) );
  AOI21_X2 U41 ( .B1(n276), .B2(n26), .A(n37), .ZN(n30) );
  INV_X4 U42 ( .A(input_base_offset), .ZN(n223) );
  INV_X4 U43 ( .A(n225), .ZN(n224) );
  INV_X4 U44 ( .A(cdf_valid), .ZN(n225) );
  AOI21_X2 U45 ( .B1(n30), .B2(reset_n), .A(n125), .ZN(n41) );
  AOI22_X2 U46 ( .A1(n277), .A2(n276), .B1(n37), .B2(input_start), .ZN(n34) );
  OAI22_X1 U47 ( .A1(n227), .A2(n196), .B1(n217), .B2(n228), .ZN(n232) );
  INV_X4 U48 ( .A(n228), .ZN(n227) );
  NAND2_X2 U49 ( .A1(n30), .A2(n31), .ZN(n25) );
  INV_X4 U50 ( .A(n25), .ZN(n275) );
  INV_X4 U51 ( .A(n26), .ZN(n229) );
  MUX2_X2 U52 ( .A(Cdf_Min[0]), .B(n217), .S(n177), .Z(n123) );
  MUX2_X2 U53 ( .A(n196), .B(Cdf_Min[0]), .S(n223), .Z(n84) );
  INV_X4 U54 ( .A(n232), .ZN(\U3/U1/Z_0 ) );
  MUX2_X2 U55 ( .A(Cdf_Min[1]), .B(n216), .S(n223), .Z(n122) );
  MUX2_X2 U56 ( .A(n201), .B(Cdf_Min[1]), .S(n223), .Z(n85) );
  MUX2_X2 U57 ( .A(n182), .B(Cdf_Min[2]), .S(n223), .Z(n86) );
  MUX2_X2 U58 ( .A(Cdf_Min[2]), .B(n214), .S(n223), .Z(n121) );
  MUX2_X2 U59 ( .A(n182), .B(n214), .S(n227), .Z(\U15/Z_2 ) );
  MUX2_X2 U60 ( .A(n183), .B(Cdf_Min[3]), .S(n177), .Z(n87) );
  MUX2_X2 U61 ( .A(Cdf_Min[3]), .B(n215), .S(n223), .Z(n120) );
  MUX2_X2 U62 ( .A(n183), .B(n215), .S(n226), .Z(\U15/Z_3 ) );
  INV_X4 U63 ( .A(\U15/Z_3 ), .ZN(n237) );
  INV_X4 U64 ( .A(n235), .ZN(n239) );
  MUX2_X2 U66 ( .A(n184), .B(Cdf_Min[4]), .S(n223), .Z(n88) );
  MUX2_X2 U67 ( .A(Cdf_Min[4]), .B(n202), .S(n223), .Z(n119) );
  MUX2_X2 U68 ( .A(n184), .B(n202), .S(n226), .Z(\U15/Z_4 ) );
  MUX2_X2 U69 ( .A(n185), .B(Cdf_Min[5]), .S(n223), .Z(n89) );
  MUX2_X2 U70 ( .A(Cdf_Min[5]), .B(n203), .S(n177), .Z(n118) );
  MUX2_X2 U73 ( .A(n185), .B(n203), .S(n227), .Z(\U15/Z_5 ) );
  NAND3_X2 U76 ( .A1(n239), .A2(n238), .A3(n237), .ZN(n240) );
  XOR2_X2 U78 ( .A(n242), .B(n218), .Z(\r312/DIFF[5] ) );
  MUX2_X2 U79 ( .A(n186), .B(Cdf_Min[6]), .S(n223), .Z(n90) );
  MUX2_X2 U80 ( .A(Cdf_Min[6]), .B(n204), .S(n223), .Z(n117) );
  MUX2_X2 U81 ( .A(n186), .B(n204), .S(n227), .Z(\U15/Z_6 ) );
  XOR2_X2 U84 ( .A(n243), .B(n241), .Z(\r312/DIFF[6] ) );
  MUX2_X2 U87 ( .A(n187), .B(Cdf_Min[7]), .S(n223), .Z(n91) );
  MUX2_X2 U90 ( .A(Cdf_Min[7]), .B(n205), .S(n177), .Z(n116) );
  MUX2_X2 U91 ( .A(n187), .B(n205), .S(n176), .Z(\U15/Z_7 ) );
  NAND3_X2 U92 ( .A1(n218), .A2(n243), .A3(n242), .ZN(n244) );
  INV_X4 U93 ( .A(n244), .ZN(n248) );
  MUX2_X2 U94 ( .A(n188), .B(Cdf_Min[8]), .S(n177), .Z(n92) );
  MUX2_X2 U95 ( .A(Cdf_Min[8]), .B(n206), .S(n177), .Z(n115) );
  MUX2_X2 U96 ( .A(n188), .B(n206), .S(n176), .Z(\U15/Z_8 ) );
  INV_X4 U97 ( .A(\U15/Z_8 ), .ZN(n247) );
  XOR2_X2 U98 ( .A(n247), .B(n245), .Z(\r312/DIFF[8] ) );
  MUX2_X2 U99 ( .A(n189), .B(Cdf_Min[9]), .S(n223), .Z(n93) );
  MUX2_X2 U100 ( .A(Cdf_Min[9]), .B(n207), .S(n223), .Z(n114) );
  MUX2_X2 U101 ( .A(n189), .B(n207), .S(n176), .Z(\U15/Z_9 ) );
  INV_X4 U102 ( .A(\U15/Z_9 ), .ZN(n251) );
  NAND3_X2 U103 ( .A1(n248), .A2(n247), .A3(n246), .ZN(n249) );
  INV_X4 U104 ( .A(n249), .ZN(n253) );
  XOR2_X2 U105 ( .A(n251), .B(n253), .Z(\r312/DIFF[9] ) );
  MUX2_X2 U106 ( .A(n190), .B(Cdf_Min[10]), .S(n223), .Z(n94) );
  MUX2_X2 U107 ( .A(Cdf_Min[10]), .B(n208), .S(n223), .Z(n113) );
  MUX2_X2 U108 ( .A(n190), .B(n208), .S(n176), .Z(\U15/Z_10 ) );
  INV_X4 U109 ( .A(\U15/Z_10 ), .ZN(n252) );
  XOR2_X2 U110 ( .A(n252), .B(n250), .Z(\r312/DIFF[10] ) );
  MUX2_X2 U111 ( .A(n191), .B(Cdf_Min[11]), .S(n223), .Z(n95) );
  MUX2_X2 U112 ( .A(Cdf_Min[11]), .B(n209), .S(n177), .Z(n112) );
  MUX2_X2 U113 ( .A(n191), .B(n209), .S(n176), .Z(\U15/Z_11 ) );
  INV_X4 U114 ( .A(\U15/Z_11 ), .ZN(n256) );
  NAND3_X2 U115 ( .A1(n253), .A2(n252), .A3(n251), .ZN(n254) );
  XOR2_X2 U116 ( .A(n256), .B(n258), .Z(\r312/DIFF[11] ) );
  MUX2_X2 U117 ( .A(n192), .B(Cdf_Min[12]), .S(n223), .Z(n96) );
  MUX2_X2 U118 ( .A(Cdf_Min[12]), .B(n210), .S(n223), .Z(n111) );
  MUX2_X2 U119 ( .A(n192), .B(n210), .S(n176), .Z(\U15/Z_12 ) );
  INV_X4 U120 ( .A(\U15/Z_12 ), .ZN(n257) );
  NAND3_X2 U121 ( .A1(n258), .A2(n257), .A3(n256), .ZN(n259) );
  MUX2_X2 U122 ( .A(n193), .B(Cdf_Min[13]), .S(n223), .Z(n97) );
  MUX2_X2 U123 ( .A(Cdf_Min[13]), .B(n211), .S(n223), .Z(n110) );
  INV_X4 U124 ( .A(n262), .ZN(n260) );
  MUX2_X2 U125 ( .A(n193), .B(n211), .S(n226), .Z(\U15/Z_13 ) );
  INV_X4 U126 ( .A(\U15/Z_13 ), .ZN(n261) );
  MUX2_X2 U127 ( .A(n194), .B(Cdf_Min[14]), .S(n177), .Z(n98) );
  MUX2_X2 U128 ( .A(Cdf_Min[14]), .B(n212), .S(n223), .Z(n109) );
  MUX2_X2 U129 ( .A(n194), .B(n212), .S(output_base_offset), .Z(\U15/Z_14 ) );
  INV_X4 U130 ( .A(\U15/Z_14 ), .ZN(n264) );
  XOR2_X2 U131 ( .A(n265), .B(n264), .Z(\r312/DIFF[14] ) );
  MUX2_X2 U132 ( .A(n195), .B(Cdf_Min[15]), .S(n223), .Z(n99) );
  MUX2_X2 U133 ( .A(Cdf_Min[15]), .B(n213), .S(n223), .Z(n108) );
  MUX2_X2 U134 ( .A(n195), .B(n213), .S(n176), .Z(\U15/Z_15 ) );
  NAND2_X2 U135 ( .A1(n265), .A2(n264), .ZN(n266) );
  NAND2_X2 U136 ( .A1(\U15/Z_15 ), .A2(n266), .ZN(n268) );
  MUX2_X2 U137 ( .A(n178), .B(Cdf_Min[16]), .S(n223), .Z(n100) );
  MUX2_X2 U138 ( .A(Cdf_Min[16]), .B(n197), .S(n177), .Z(n107) );
  MUX2_X2 U139 ( .A(n178), .B(n197), .S(output_base_offset), .Z(\U15/Z_16 ) );
  INV_X4 U140 ( .A(\U15/Z_16 ), .ZN(n267) );
  XOR2_X2 U141 ( .A(n268), .B(n267), .Z(\r312/DIFF[16] ) );
  MUX2_X2 U142 ( .A(n179), .B(Cdf_Min[17]), .S(n223), .Z(n101) );
  MUX2_X2 U143 ( .A(Cdf_Min[17]), .B(n198), .S(n223), .Z(n106) );
  MUX2_X2 U144 ( .A(n179), .B(n198), .S(n176), .Z(\U15/Z_17 ) );
  INV_X4 U145 ( .A(\U15/Z_17 ), .ZN(n270) );
  NAND2_X2 U146 ( .A1(n268), .A2(n267), .ZN(n269) );
  INV_X4 U147 ( .A(n269), .ZN(n271) );
  XOR2_X2 U148 ( .A(n270), .B(n271), .Z(\r312/DIFF[17] ) );
  MUX2_X2 U149 ( .A(n180), .B(Cdf_Min[18]), .S(n223), .Z(n102) );
  MUX2_X2 U150 ( .A(Cdf_Min[18]), .B(n199), .S(n223), .Z(n105) );
  NAND2_X2 U151 ( .A1(n271), .A2(n270), .ZN(n272) );
  MUX2_X2 U152 ( .A(n180), .B(n199), .S(output_base_offset), .Z(\U15/Z_18 ) );
  MUX2_X2 U153 ( .A(n181), .B(Cdf_Min[19]), .S(n223), .Z(n103) );
  MUX2_X2 U154 ( .A(Cdf_Min[19]), .B(n200), .S(n223), .Z(n104) );
  NAND2_X2 U155 ( .A1(\U15/Z_18 ), .A2(n272), .ZN(n273) );
  MUX2_X2 U156 ( .A(n181), .B(n200), .S(n176), .Z(\U15/Z_19 ) );
  INV_X4 U157 ( .A(n41), .ZN(n274) );
  INV_X4 U158 ( .A(\U10/DATA2_0 ), .ZN(n276) );
  INV_X4 U159 ( .A(n37), .ZN(n278) );
  INV_X4 U160 ( .A(n31), .ZN(n279) );
endmodule


module input_pipeline ( start, clock, rst_n, m1ReadBus, m2ReadBus, 
        inputBaseOffset, m1ReadAddr, m2ReadAddr, m2WriteAddr, m3WriteAddr, 
        m2WriteBus, m3WriteBus, m2WE, m3WE, input_done );
  input [127:0] m1ReadBus;
  input [35:0] m2ReadBus;
  output [15:0] m1ReadAddr;
  output [15:0] m2ReadAddr;
  output [15:0] m2WriteAddr;
  output [15:0] m3WriteAddr;
  output [127:0] m2WriteBus;
  output [127:0] m3WriteBus;
  input start, clock, rst_n, inputBaseOffset;
  output m2WE, m3WE, input_done;
  wire   n448, n501, \U3/U1/Z_0 , \U3/U1/DATA2_0 , \U3/U1/DATA2_1 ,
         \U3/U1/DATA2_2 , \U3/U1/DATA2_3 , \U3/U1/DATA2_4 , \U3/U1/DATA2_5 ,
         \U3/U1/DATA2_6 , \U3/U1/DATA2_7 , \U3/U1/DATA2_8 , \U3/U1/DATA2_9 ,
         \U3/U1/DATA2_10 , \U3/U1/DATA2_11 , \U3/U1/DATA2_12 ,
         \U3/U1/DATA2_13 , \U3/U1/DATA2_14 , \U3/U1/DATA2_15 ,
         \U3/U1/DATA2_16 , \U3/U1/DATA2_17 , \U3/U1/DATA2_18 ,
         \U3/U1/DATA2_19 , \U3/U1/DATA2_20 , \U3/U1/DATA2_21 ,
         \U3/U1/DATA2_22 , \U3/U1/DATA2_23 , \U3/U1/DATA2_24 ,
         \U3/U1/DATA2_25 , \U3/U1/DATA2_26 , \U3/U1/DATA2_27 ,
         \U3/U1/DATA2_28 , \U3/U1/DATA2_29 , \U3/U1/DATA2_30 ,
         \U3/U1/DATA2_31 , \U3/U1/DATA2_32 , \U3/U1/DATA2_33 ,
         \U3/U1/DATA2_34 , \U3/U1/DATA2_35 , \U3/U1/DATA1_0 , \U3/U1/DATA1_1 ,
         \U3/U1/DATA1_2 , \U3/U1/DATA1_3 , \U3/U1/DATA1_4 , \U3/U1/DATA1_5 ,
         \U3/U1/DATA1_6 , \U3/U1/DATA1_7 , \U3/U1/DATA1_8 , \U3/U1/DATA1_9 ,
         \U3/U1/DATA1_10 , \U3/U1/DATA1_11 , \U3/U1/DATA1_12 ,
         \U3/U1/DATA1_13 , \U3/U1/DATA1_14 , \U3/U1/DATA1_15 ,
         \U3/U1/DATA1_16 , \U3/U1/DATA1_17 , \U3/U1/DATA1_18 ,
         \U3/U1/DATA1_19 , \U3/U1/DATA1_20 , \U3/U1/DATA1_21 ,
         \U3/U1/DATA1_22 , \U3/U1/DATA1_23 , \U3/U1/DATA1_24 ,
         \U3/U1/DATA1_25 , \U3/U1/DATA1_26 , \U3/U1/DATA1_27 ,
         \U3/U1/DATA1_28 , \U3/U1/DATA1_29 , \U3/U1/DATA1_30 ,
         \U3/U1/DATA1_31 , \U3/U1/DATA1_32 , \U3/U1/DATA1_33 ,
         \U3/U1/DATA1_34 , \U3/U1/DATA1_35 , \U35/DATA2_0 , \U35/DATA2_1 ,
         \U35/DATA2_2 , \U35/DATA2_3 , \U35/DATA2_4 , \U35/DATA2_5 ,
         \U35/DATA2_6 , \U35/DATA2_7 , \U35/DATA2_8 , \U35/DATA2_9 ,
         \U35/DATA2_10 , \U35/DATA2_11 , \U35/DATA2_12 , \U35/DATA2_13 ,
         \U35/DATA2_14 , \U35/DATA2_15 , \U35/DATA2_16 , \U35/DATA2_17 ,
         \U35/DATA2_18 , \U35/DATA2_19 , \U35/DATA2_20 , \U35/DATA2_21 ,
         \U35/DATA2_22 , \U35/DATA2_23 , \U35/DATA2_24 , \U35/DATA2_25 ,
         \U35/DATA2_26 , \U35/DATA2_27 , \U35/DATA2_28 , \U35/DATA2_29 ,
         \U35/DATA2_30 , \U35/DATA2_31 , \U35/DATA2_32 , \U35/DATA2_33 ,
         \U35/DATA2_34 , \U35/DATA2_35 , \U35/DATA2_36 , \U35/DATA2_37 ,
         \U35/DATA2_38 , \U35/DATA2_39 , \U35/DATA2_40 , \U35/DATA2_41 ,
         \U35/DATA2_42 , \U35/DATA2_43 , \U35/DATA2_44 , \U35/DATA2_45 ,
         \U35/DATA2_46 , \U35/DATA2_47 , \U35/DATA2_48 , \U35/DATA2_49 ,
         \U35/DATA2_50 , \U35/DATA2_51 , \U35/DATA2_52 , \U35/DATA2_53 ,
         \U35/DATA2_54 , \U35/DATA2_55 , \U35/DATA2_56 , \U35/DATA2_57 ,
         \U35/DATA2_58 , \U35/DATA2_59 , \U35/DATA2_60 , \U35/DATA2_61 ,
         \U35/DATA2_62 , \U35/DATA2_63 , \U35/DATA2_64 , \U35/DATA2_65 ,
         \U35/DATA2_66 , \U35/DATA2_67 , \U35/DATA2_68 , \U35/DATA2_69 ,
         \U35/DATA2_70 , \U35/DATA1_7 , \U35/DATA1_8 , \U35/DATA1_9 ,
         \U35/DATA1_10 , \U35/DATA1_11 , \U35/DATA1_12 , \U35/DATA1_13 ,
         \U35/DATA1_14 , \U35/DATA1_15 , \U35/DATA1_16 , \U35/DATA1_17 ,
         \U35/DATA1_18 , \U35/DATA1_19 , \U35/DATA1_20 , \U35/DATA1_21 ,
         \U35/DATA1_22 , \U35/DATA1_23 , \U35/DATA1_24 , \U35/DATA1_25 ,
         \U35/DATA1_26 , \U35/DATA1_27 , \U35/DATA1_28 , \U35/DATA1_29 ,
         \U35/DATA1_30 , \U35/DATA1_31 , \U35/DATA1_32 , \U35/DATA1_33 ,
         \U35/DATA1_34 , \U35/DATA1_35 , \U35/DATA1_36 , \U35/DATA1_37 ,
         \U35/DATA1_38 , \U35/DATA1_39 , \U35/DATA1_40 , \U35/DATA1_41 ,
         \U35/DATA1_42 , \U35/DATA1_43 , \U35/DATA1_44 , \U35/DATA1_45 ,
         \U35/DATA1_46 , \U35/DATA1_47 , \U35/DATA1_48 , \U35/DATA1_49 ,
         \U35/DATA1_50 , \U35/DATA1_51 , \U35/DATA1_52 , \U35/DATA1_53 ,
         \U35/DATA1_54 , \U35/DATA1_55 , \U35/DATA1_56 , \U35/DATA1_57 ,
         \U35/DATA1_58 , \U35/DATA1_59 , \U35/DATA1_60 , \U35/DATA1_61 ,
         \U35/DATA1_62 , \U35/DATA1_63 , \U28/DATA2_0 , \U28/DATA2_1 ,
         \U28/DATA2_2 , \U28/DATA2_3 , \U28/DATA2_4 , \U28/DATA2_5 ,
         \U28/DATA2_6 , \U28/DATA2_7 , \U28/DATA2_8 , \U28/DATA2_9 ,
         \U28/DATA2_10 , \U28/DATA2_11 , \U28/DATA2_12 , \U28/DATA2_13 ,
         \U28/DATA2_14 , \U28/DATA2_15 , \U28/DATA2_16 , \U28/DATA2_17 ,
         \U28/DATA2_18 , \U28/DATA2_19 , \U28/DATA2_20 , \U28/DATA2_21 ,
         \U28/DATA2_22 , \U28/DATA2_23 , \U28/DATA2_24 , \U28/DATA2_25 ,
         \U28/DATA2_26 , \U28/DATA2_27 , \U28/DATA2_28 , \U28/DATA2_29 ,
         \U28/DATA2_30 , \U28/DATA2_31 , \U28/DATA2_32 , \U28/DATA2_33 ,
         \U28/DATA2_34 , \U28/DATA2_35 , \U28/DATA1_0 , \U28/DATA1_1 ,
         \U28/DATA1_2 , \U28/DATA1_3 , \U28/DATA1_4 , \U28/DATA1_5 ,
         \U28/DATA1_6 , \U28/DATA1_7 , \U28/DATA1_8 , \U28/DATA1_9 ,
         \U28/DATA1_10 , \U28/DATA1_11 , \U28/DATA1_12 , \U28/DATA1_13 ,
         \U28/DATA1_14 , \U28/DATA1_15 , \U28/DATA1_16 , \U28/DATA1_17 ,
         \U28/DATA1_18 , \U28/DATA1_19 , \U28/DATA1_20 , \U28/DATA1_21 ,
         \U28/DATA1_22 , \U28/DATA1_23 , \U28/DATA1_24 , \U28/DATA1_25 ,
         \U28/DATA1_26 , \U28/DATA1_27 , \U28/DATA1_28 , \U28/DATA1_29 ,
         \U28/DATA1_30 , \U28/DATA1_31 , \U28/DATA1_32 , \U28/DATA1_33 ,
         \U28/DATA1_34 , \U28/DATA1_35 , \U26/Z_0 , \U26/DATA1_0 , \U25/Z_0 ,
         \U25/DATA1_0 , \U23/Z_0 , \U23/DATA1_0 , \U22/Z_0 , \U22/DATA1_0 ,
         \U21/Z_0 , \U21/Z_1 , \U21/Z_2 , \U21/Z_3 , \U21/Z_4 , \U21/Z_5 ,
         \U21/Z_6 , \U21/Z_7 , \U21/DATA1_0 , \U21/DATA1_1 , \U21/DATA1_2 ,
         \U21/DATA1_3 , \U21/DATA1_4 , \U21/DATA1_5 , \U21/DATA1_6 ,
         \U21/DATA1_7 , \U20/Z_0 , \U20/Z_1 , \U20/Z_2 , \U20/Z_3 , \U20/Z_4 ,
         \U20/Z_5 , \U20/Z_6 , \U20/Z_7 , \U20/Z_8 , \U20/Z_9 , \U20/Z_10 ,
         \U20/Z_11 , \U20/Z_12 , \U20/Z_13 , \U20/Z_14 , \U20/Z_15 ,
         \U20/Z_16 , \U20/Z_17 , \U20/Z_18 , \U20/Z_19 , \U20/Z_20 ,
         \U20/Z_21 , \U20/Z_22 , \U20/Z_23 , \U20/Z_24 , \U20/Z_25 ,
         \U20/Z_26 , \U20/Z_27 , \U20/Z_28 , \U20/Z_29 , \U20/Z_30 ,
         \U20/Z_31 , \U20/Z_32 , \U20/Z_33 , \U20/Z_34 , \U20/Z_35 , \U19/Z_0 ,
         \U19/DATA1_0 , \U18/Z_0 , \U18/DATA1_0 , \U17/Z_0 , \U17/Z_1 ,
         \U17/Z_2 , \U17/Z_3 , \U17/Z_4 , \U17/Z_5 , \U17/Z_6 , \U17/Z_7 ,
         \U17/DATA1_2 , \U17/DATA1_6 , \U17/DATA1_7 , \U16/Z_1 , \U16/Z_2 ,
         \U16/Z_3 , \U16/Z_4 , \U16/Z_5 , \U16/Z_6 , \U16/Z_7 , \U16/Z_8 ,
         \U16/Z_9 , \U16/Z_10 , \U16/Z_11 , \U16/Z_12 , \U16/Z_13 , \U16/Z_14 ,
         \U16/Z_15 , \U16/Z_16 , \U16/Z_17 , \U16/Z_18 , \U16/Z_19 ,
         \U16/Z_20 , \U16/Z_22 , \U16/Z_24 , \U16/Z_26 , \U16/Z_28 ,
         \U16/Z_30 , \U16/Z_32 , \U16/Z_34 , \U16/Z_35 , \U16/DATA1_21 ,
         \U16/DATA1_23 , \U16/DATA1_25 , \U16/DATA1_27 , \U16/DATA1_29 ,
         \U16/DATA1_31 , \U16/DATA1_33 , \U15/DATA1_3 , \U15/DATA1_4 ,
         \U15/DATA1_5 , \U15/DATA1_6 , \U14/Z_0 , \U5/DATA1_0 , \U5/DATA1_1 ,
         \U5/DATA1_2 , \U5/DATA1_3 , \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 ,
         \U5/DATA1_7 , \U5/DATA1_8 , \U5/DATA1_9 , \U5/DATA1_10 ,
         \U5/DATA1_11 , \U5/DATA1_12 , \U5/DATA1_13 , \U5/DATA1_14 ,
         \U5/DATA1_15 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 , \eq_122/B[7] ,
         \eq_122/B[6] , \eq_122/B[5] , \eq_122/B[4] , \eq_122/B[3] ,
         \eq_122/B[2] , \eq_122/B[1] , \eq_122/B[0] , \eq_62/B[7] ,
         \eq_62/B[6] , \eq_62/B[5] , \eq_62/B[4] , \eq_62/B[3] , \eq_62/B[2] ,
         \eq_62/B[1] , \eq_62/B[0] , n20, n21, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n113, n115, n121, n123, n127, n128, n147, n148, n149, n190, n191,
         n192, n201, n205, n207, n208, n212, n213, n214, n218, n219, n220,
         n225, n227, n230, n233, n236, n237, n238, n239, n240, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n319, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n370, n371, n372, n373, n420, n421, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;
  assign \U35/DATA2_0  = m1ReadBus[0];
  assign \U35/DATA2_1  = m1ReadBus[1];
  assign \U35/DATA2_2  = m1ReadBus[2];
  assign \U35/DATA2_3  = m1ReadBus[3];
  assign \U35/DATA2_4  = m1ReadBus[4];
  assign \U35/DATA2_5  = m1ReadBus[5];
  assign \U35/DATA2_6  = m1ReadBus[6];
  assign \U35/DATA2_7  = m1ReadBus[7];
  assign \U35/DATA2_8  = m1ReadBus[8];
  assign \U35/DATA2_9  = m1ReadBus[9];
  assign \U35/DATA2_10  = m1ReadBus[10];
  assign \U35/DATA2_11  = m1ReadBus[11];
  assign \U35/DATA2_12  = m1ReadBus[12];
  assign \U35/DATA2_13  = m1ReadBus[13];
  assign \U35/DATA2_14  = m1ReadBus[14];
  assign \U35/DATA2_15  = m1ReadBus[15];
  assign \U35/DATA2_16  = m1ReadBus[16];
  assign \U35/DATA2_17  = m1ReadBus[17];
  assign \U35/DATA2_18  = m1ReadBus[18];
  assign \U35/DATA2_19  = m1ReadBus[19];
  assign \U35/DATA2_20  = m1ReadBus[20];
  assign \U35/DATA2_21  = m1ReadBus[21];
  assign \U35/DATA2_22  = m1ReadBus[22];
  assign \U35/DATA2_23  = m1ReadBus[23];
  assign \U35/DATA2_24  = m1ReadBus[24];
  assign \U35/DATA2_25  = m1ReadBus[25];
  assign \U35/DATA2_26  = m1ReadBus[26];
  assign \U35/DATA2_27  = m1ReadBus[27];
  assign \U35/DATA2_28  = m1ReadBus[28];
  assign \U35/DATA2_29  = m1ReadBus[29];
  assign \U35/DATA2_30  = m1ReadBus[30];
  assign \U35/DATA2_31  = m1ReadBus[31];
  assign \U35/DATA2_32  = m1ReadBus[32];
  assign \U35/DATA2_33  = m1ReadBus[33];
  assign \U35/DATA2_34  = m1ReadBus[34];
  assign \U35/DATA2_35  = m1ReadBus[35];
  assign \U35/DATA2_36  = m1ReadBus[36];
  assign \U35/DATA2_37  = m1ReadBus[37];
  assign \U35/DATA2_38  = m1ReadBus[38];
  assign \U35/DATA2_39  = m1ReadBus[39];
  assign \U35/DATA2_40  = m1ReadBus[40];
  assign \U35/DATA2_41  = m1ReadBus[41];
  assign \U35/DATA2_42  = m1ReadBus[42];
  assign \U35/DATA2_43  = m1ReadBus[43];
  assign \U35/DATA2_44  = m1ReadBus[44];
  assign \U35/DATA2_45  = m1ReadBus[45];
  assign \U35/DATA2_46  = m1ReadBus[46];
  assign \U35/DATA2_47  = m1ReadBus[47];
  assign \U35/DATA2_48  = m1ReadBus[48];
  assign \U35/DATA2_49  = m1ReadBus[49];
  assign \U35/DATA2_50  = m1ReadBus[50];
  assign \U35/DATA2_51  = m1ReadBus[51];
  assign \U35/DATA2_52  = m1ReadBus[52];
  assign \U35/DATA2_53  = m1ReadBus[53];
  assign \U35/DATA2_54  = m1ReadBus[54];
  assign \U35/DATA2_55  = m1ReadBus[55];
  assign \U35/DATA2_56  = m1ReadBus[56];
  assign \U35/DATA2_57  = m1ReadBus[57];
  assign \U35/DATA2_58  = m1ReadBus[58];
  assign \U35/DATA2_59  = m1ReadBus[59];
  assign \U35/DATA2_60  = m1ReadBus[60];
  assign \U35/DATA2_61  = m1ReadBus[61];
  assign \U35/DATA2_62  = m1ReadBus[62];
  assign \U35/DATA2_63  = m1ReadBus[63];
  assign \U35/DATA2_64  = m1ReadBus[64];
  assign \U35/DATA2_65  = m1ReadBus[65];
  assign \U35/DATA2_66  = m1ReadBus[66];
  assign \U35/DATA2_67  = m1ReadBus[67];
  assign \U35/DATA2_68  = m1ReadBus[68];
  assign \U35/DATA2_69  = m1ReadBus[69];
  assign \U35/DATA2_70  = m1ReadBus[70];
  assign \U35/DATA1_7  = m1ReadBus[71];
  assign \U35/DATA1_8  = m1ReadBus[72];
  assign \U35/DATA1_9  = m1ReadBus[73];
  assign \U35/DATA1_10  = m1ReadBus[74];
  assign \U35/DATA1_11  = m1ReadBus[75];
  assign \U35/DATA1_12  = m1ReadBus[76];
  assign \U35/DATA1_13  = m1ReadBus[77];
  assign \U35/DATA1_14  = m1ReadBus[78];
  assign \U35/DATA1_15  = m1ReadBus[79];
  assign \U35/DATA1_16  = m1ReadBus[80];
  assign \U35/DATA1_17  = m1ReadBus[81];
  assign \U35/DATA1_18  = m1ReadBus[82];
  assign \U35/DATA1_19  = m1ReadBus[83];
  assign \U35/DATA1_20  = m1ReadBus[84];
  assign \U35/DATA1_21  = m1ReadBus[85];
  assign \U35/DATA1_22  = m1ReadBus[86];
  assign \U35/DATA1_23  = m1ReadBus[87];
  assign \U35/DATA1_24  = m1ReadBus[88];
  assign \U35/DATA1_25  = m1ReadBus[89];
  assign \U35/DATA1_26  = m1ReadBus[90];
  assign \U35/DATA1_27  = m1ReadBus[91];
  assign \U35/DATA1_28  = m1ReadBus[92];
  assign \U35/DATA1_29  = m1ReadBus[93];
  assign \U35/DATA1_30  = m1ReadBus[94];
  assign \U35/DATA1_31  = m1ReadBus[95];
  assign \U35/DATA1_32  = m1ReadBus[96];
  assign \U35/DATA1_33  = m1ReadBus[97];
  assign \U35/DATA1_34  = m1ReadBus[98];
  assign \U35/DATA1_35  = m1ReadBus[99];
  assign \U35/DATA1_36  = m1ReadBus[100];
  assign \U35/DATA1_37  = m1ReadBus[101];
  assign \U35/DATA1_38  = m1ReadBus[102];
  assign \U35/DATA1_39  = m1ReadBus[103];
  assign \U35/DATA1_40  = m1ReadBus[104];
  assign \U35/DATA1_41  = m1ReadBus[105];
  assign \U35/DATA1_42  = m1ReadBus[106];
  assign \U35/DATA1_43  = m1ReadBus[107];
  assign \U35/DATA1_44  = m1ReadBus[108];
  assign \U35/DATA1_45  = m1ReadBus[109];
  assign \U35/DATA1_46  = m1ReadBus[110];
  assign \U35/DATA1_47  = m1ReadBus[111];
  assign \U35/DATA1_48  = m1ReadBus[112];
  assign \U35/DATA1_49  = m1ReadBus[113];
  assign \U35/DATA1_50  = m1ReadBus[114];
  assign \U35/DATA1_51  = m1ReadBus[115];
  assign \U35/DATA1_52  = m1ReadBus[116];
  assign \U35/DATA1_53  = m1ReadBus[117];
  assign \U35/DATA1_54  = m1ReadBus[118];
  assign \U35/DATA1_55  = m1ReadBus[119];
  assign \U35/DATA1_56  = m1ReadBus[120];
  assign \U35/DATA1_57  = m1ReadBus[121];
  assign \U35/DATA1_58  = m1ReadBus[122];
  assign \U35/DATA1_59  = m1ReadBus[123];
  assign \U35/DATA1_60  = m1ReadBus[124];
  assign \U35/DATA1_61  = m1ReadBus[125];
  assign \U35/DATA1_62  = m1ReadBus[126];
  assign \U35/DATA1_63  = m1ReadBus[127];
  assign \U28/DATA2_0  = m2ReadBus[0];
  assign \U28/DATA2_1  = m2ReadBus[1];
  assign \U28/DATA2_2  = m2ReadBus[2];
  assign \U28/DATA2_3  = m2ReadBus[3];
  assign \U28/DATA2_4  = m2ReadBus[4];
  assign \U28/DATA2_5  = m2ReadBus[5];
  assign \U28/DATA2_6  = m2ReadBus[6];
  assign \U28/DATA2_7  = m2ReadBus[7];
  assign \U28/DATA2_8  = m2ReadBus[8];
  assign \U28/DATA2_9  = m2ReadBus[9];
  assign \U28/DATA2_10  = m2ReadBus[10];
  assign \U28/DATA2_11  = m2ReadBus[11];
  assign \U28/DATA2_12  = m2ReadBus[12];
  assign \U28/DATA2_13  = m2ReadBus[13];
  assign \U28/DATA2_14  = m2ReadBus[14];
  assign \U28/DATA2_15  = m2ReadBus[15];
  assign \U28/DATA2_16  = m2ReadBus[16];
  assign \U28/DATA2_17  = m2ReadBus[17];
  assign \U28/DATA2_18  = m2ReadBus[18];
  assign \U28/DATA2_19  = m2ReadBus[19];
  assign \U28/DATA2_20  = m2ReadBus[20];
  assign \U28/DATA2_21  = m2ReadBus[21];
  assign \U28/DATA2_22  = m2ReadBus[22];
  assign \U28/DATA2_23  = m2ReadBus[23];
  assign \U28/DATA2_24  = m2ReadBus[24];
  assign \U28/DATA2_25  = m2ReadBus[25];
  assign \U28/DATA2_26  = m2ReadBus[26];
  assign \U28/DATA2_27  = m2ReadBus[27];
  assign \U28/DATA2_28  = m2ReadBus[28];
  assign \U28/DATA2_29  = m2ReadBus[29];
  assign \U28/DATA2_30  = m2ReadBus[30];
  assign \U28/DATA2_31  = m2ReadBus[31];
  assign \U28/DATA2_32  = m2ReadBus[32];
  assign \U28/DATA2_33  = m2ReadBus[33];
  assign \U28/DATA2_34  = m2ReadBus[34];
  assign \U28/DATA2_35  = m2ReadBus[35];
  assign m2WriteBus[0] = \U28/DATA1_0 ;
  assign m2WriteBus[1] = \U28/DATA1_1 ;
  assign m2WriteBus[2] = \U28/DATA1_2 ;
  assign m2WriteBus[3] = \U28/DATA1_3 ;
  assign m2WriteBus[4] = \U28/DATA1_4 ;
  assign m2WriteBus[5] = \U28/DATA1_5 ;
  assign m2WriteBus[6] = \U28/DATA1_6 ;
  assign m2WriteBus[7] = \U28/DATA1_7 ;
  assign m2WriteBus[8] = \U28/DATA1_8 ;
  assign m2WriteBus[9] = \U28/DATA1_9 ;
  assign m2WriteBus[10] = \U28/DATA1_10 ;
  assign m2WriteBus[11] = \U28/DATA1_11 ;
  assign m2WriteBus[12] = \U28/DATA1_12 ;
  assign m2WriteBus[13] = \U28/DATA1_13 ;
  assign m2WriteBus[14] = \U28/DATA1_14 ;
  assign m2WriteBus[15] = \U28/DATA1_15 ;
  assign m2WriteBus[16] = \U28/DATA1_16 ;
  assign m2WriteBus[17] = \U28/DATA1_17 ;
  assign m2WriteBus[18] = \U28/DATA1_18 ;
  assign m2WriteBus[19] = \U28/DATA1_19 ;
  assign m2WriteBus[20] = \U28/DATA1_20 ;
  assign m2WriteBus[21] = \U28/DATA1_21 ;
  assign m2WriteBus[22] = \U28/DATA1_22 ;
  assign m2WriteBus[23] = \U28/DATA1_23 ;
  assign m2WriteBus[24] = \U28/DATA1_24 ;
  assign m2WriteBus[25] = \U28/DATA1_25 ;
  assign m2WriteBus[26] = \U28/DATA1_26 ;
  assign m2WriteBus[27] = \U28/DATA1_27 ;
  assign m2WriteBus[28] = \U28/DATA1_28 ;
  assign m2WriteBus[29] = \U28/DATA1_29 ;
  assign m2WriteBus[30] = \U28/DATA1_30 ;
  assign m2WriteBus[31] = \U28/DATA1_31 ;
  assign m2WriteBus[32] = \U28/DATA1_32 ;
  assign m2WriteBus[33] = \U28/DATA1_33 ;
  assign m2WriteBus[34] = \U28/DATA1_34 ;
  assign m2WriteBus[35] = \U28/DATA1_35 ;
  assign m2ReadAddr[0] = \U21/DATA1_0 ;
  assign m2ReadAddr[1] = \U21/DATA1_1 ;
  assign m2ReadAddr[2] = \U21/DATA1_2 ;
  assign m2ReadAddr[3] = \U21/DATA1_3 ;
  assign m2ReadAddr[4] = \U21/DATA1_4 ;
  assign m2ReadAddr[5] = \U21/DATA1_5 ;
  assign m2ReadAddr[6] = \U21/DATA1_6 ;
  assign m2ReadAddr[7] = \U21/DATA1_7 ;
  assign m1ReadAddr[0] = \U5/DATA1_0 ;
  assign m1ReadAddr[1] = \U5/DATA1_1 ;
  assign m1ReadAddr[2] = \U5/DATA1_2 ;
  assign m1ReadAddr[3] = \U5/DATA1_3 ;
  assign m1ReadAddr[4] = \U5/DATA1_4 ;
  assign m1ReadAddr[5] = \U5/DATA1_5 ;
  assign m1ReadAddr[6] = \U5/DATA1_6 ;
  assign m1ReadAddr[7] = \U5/DATA1_7 ;
  assign m1ReadAddr[8] = \U5/DATA1_8 ;
  assign m1ReadAddr[9] = \U5/DATA1_9 ;
  assign m1ReadAddr[10] = \U5/DATA1_10 ;
  assign m1ReadAddr[11] = \U5/DATA1_11 ;
  assign m1ReadAddr[12] = \U5/DATA1_12 ;
  assign m1ReadAddr[13] = \U5/DATA1_13 ;
  assign m1ReadAddr[14] = \U5/DATA1_14 ;
  assign m1ReadAddr[15] = \U5/DATA1_15 ;
  assign m2WriteAddr[7] = \eq_62/B[7] ;
  assign m2WriteAddr[6] = \eq_62/B[6] ;
  assign m2WriteAddr[5] = \eq_62/B[5] ;
  assign m2WriteAddr[4] = \eq_62/B[4] ;
  assign m2WriteAddr[3] = \eq_62/B[3] ;
  assign m2WriteAddr[2] = \eq_62/B[2] ;
  assign m2WriteAddr[1] = \eq_62/B[1] ;
  assign m2WriteAddr[0] = \eq_62/B[0] ;

  SDFFR_X2 write_enable_reg ( .D(1'b1), .SI(n148), .SE(n1460), .CK(clock), 
        .RN(rst_n), .Q(\U25/DATA1_0 ) );
  DFFR_X1 m2WE_Accum_reg ( .D(\U18/Z_0 ), .CK(clock), .RN(n1529), .Q(n501), 
        .QN(n20) );
  DFFR_X1 done_enable_reg ( .D(n1806), .CK(clock), .RN(n1529), .Q(
        \U26/DATA1_0 ) );
  DFFR_X1 \pipelineCounter_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n1529), .Q(
        \U15/DATA1_5 ), .QN(n115) );
  DFFR_X1 \pipelineCounter_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n1529), .Q(
        \U15/DATA1_6 ), .QN(n113) );
  DFFR_X1 \readInitial_FS_reg[7]  ( .D(\U21/Z_7 ), .CK(clock), .RN(n1531), .Q(
        \U17/DATA1_7 ), .QN(n1472) );
  DFFR_X1 \readInitial_Accum_reg[7]  ( .D(\U17/Z_7 ), .CK(clock), .RN(n1531), 
        .Q(\eq_122/B[7] ) );
  SDFFR_X2 \readInitial_FI_reg[6]  ( .D(n1521), .SI(1'b0), .SE(n218), .CK(
        clock), .RN(rst_n), .Q(\U21/DATA1_6 ), .QN(n1545) );
  DFFR_X1 \readInitial_Accum_reg[6]  ( .D(\U17/Z_6 ), .CK(clock), .RN(n1531), 
        .Q(\eq_122/B[6] ) );
  SDFFR_X2 \readInitial_FI_reg[5]  ( .D(n1521), .SI(1'b0), .SE(n1809), .CK(
        clock), .RN(rst_n), .Q(\U21/DATA1_5 ), .QN(n1541) );
  SDFFR_X2 \readInitial_FI_reg[4]  ( .D(n1521), .SI(1'b0), .SE(n230), .CK(
        clock), .RN(rst_n), .Q(\U21/DATA1_4 ), .QN(n1543) );
  SDFFR_X2 \readInitial_FI_reg[3]  ( .D(n1521), .SI(1'b0), .SE(n294), .CK(
        clock), .RN(rst_n), .Q(\U21/DATA1_3 ), .QN(n1544) );
  SDFFR_X2 \readInitial_FI_reg[2]  ( .D(n1521), .SI(1'b0), .SE(n236), .CK(
        clock), .RN(rst_n), .Q(\U21/DATA1_2 ), .QN(n1538) );
  DFFR_X1 \readInitial_FS_reg[2]  ( .D(\U21/Z_2 ), .CK(clock), .RN(n1532), .Q(
        \U17/DATA1_2 ), .QN(n1462) );
  DFFR_X1 \readInitial_Accum_reg[2]  ( .D(\U17/Z_2 ), .CK(clock), .RN(n1532), 
        .Q(\eq_122/B[2] ) );
  SDFFR_X2 \readInitial_FI_reg[1]  ( .D(n1521), .SI(1'b0), .SE(n1808), .CK(
        clock), .RN(rst_n), .Q(\U21/DATA1_1 ), .QN(n1539) );
  DFFR_X1 \readInitial_FS_reg[1]  ( .D(\U21/Z_1 ), .CK(clock), .RN(n1532), 
        .QN(n1458) );
  SDFFR_X2 \readInitial_FI_reg[0]  ( .D(n1521), .SI(1'b0), .SE(n1810), .CK(
        clock), .RN(rst_n), .Q(\U21/DATA1_0 ), .QN(n1546) );
  DFFR_X1 \readInitial_FS_reg[0]  ( .D(\U21/Z_0 ), .CK(clock), .RN(n1532), 
        .QN(n1457) );
  DFFR_X1 \scratchVal_FS_reg[0]  ( .D(\U20/Z_0 ), .CK(clock), .RN(n1532), .Q(
        \U3/U1/DATA2_0 ) );
  DFFR_X1 \scratchVal_Accum_reg[1]  ( .D(\U16/Z_1 ), .CK(clock), .RN(n1532), 
        .Q(\U3/U1/DATA1_1 ), .QN(n56) );
  DFFR_X1 \scratchVal_Accum_reg[2]  ( .D(\U16/Z_2 ), .CK(clock), .RN(n1532), 
        .Q(\U3/U1/DATA1_2 ), .QN(n55) );
  DFFR_X1 \scratchVal_Accum_reg[3]  ( .D(\U16/Z_3 ), .CK(clock), .RN(n1532), 
        .Q(\U3/U1/DATA1_3 ), .QN(n54) );
  DFFR_X1 \scratchVal_Accum_reg[4]  ( .D(\U16/Z_4 ), .CK(clock), .RN(n1532), 
        .Q(\U3/U1/DATA1_4 ), .QN(n53) );
  DFFR_X1 \scratchVal_Accum_reg[5]  ( .D(\U16/Z_5 ), .CK(clock), .RN(n1532), 
        .Q(\U3/U1/DATA1_5 ), .QN(n52) );
  DFFR_X1 \scratchVal_Accum_reg[6]  ( .D(\U16/Z_6 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_6 ), .QN(n51) );
  DFFR_X1 \scratchVal_Accum_reg[7]  ( .D(\U16/Z_7 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_7 ), .QN(n50) );
  DFFR_X1 \scratchVal_Accum_reg[8]  ( .D(\U16/Z_8 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_8 ), .QN(n49) );
  DFFR_X1 \scratchVal_Accum_reg[9]  ( .D(\U16/Z_9 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_9 ), .QN(n48) );
  DFFR_X1 \scratchVal_Accum_reg[10]  ( .D(\U16/Z_10 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_10 ), .QN(n47) );
  DFFR_X1 \scratchVal_Accum_reg[11]  ( .D(\U16/Z_11 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_11 ), .QN(n46) );
  DFFR_X1 \scratchVal_Accum_reg[12]  ( .D(\U16/Z_12 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_12 ), .QN(n45) );
  DFFR_X1 \scratchVal_Accum_reg[13]  ( .D(\U16/Z_13 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_13 ), .QN(n44) );
  DFFR_X1 \scratchVal_Accum_reg[14]  ( .D(\U16/Z_14 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_14 ), .QN(n42) );
  DFFR_X1 \scratchVal_Accum_reg[15]  ( .D(\U16/Z_15 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_15 ), .QN(n41) );
  DFFR_X1 \scratchVal_Accum_reg[17]  ( .D(\U16/Z_17 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA1_17 ), .QN(n39) );
  DFFR_X1 \scratchVal_Accum_reg[18]  ( .D(\U16/Z_18 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_18 ), .QN(n38) );
  DFFR_X1 \scratchVal_Accum_reg[19]  ( .D(\U16/Z_19 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA1_19 ), .QN(n37) );
  DFFR_X1 \scratchVal_Accum_reg[20]  ( .D(\U16/Z_20 ), .CK(clock), .RN(n1529), 
        .Q(\U3/U1/DATA1_20 ), .QN(n36) );
  DFFR_X1 \scratchVal_FS_reg[20]  ( .D(\U20/Z_20 ), .CK(clock), .RN(n1529), 
        .Q(\U3/U1/DATA2_20 ) );
  DFFS_X2 \scratchVal_FS_reg[21]  ( .D(\U20/Z_21 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA2_21 ) );
  DFFR_X1 \scratchVal_Accum_reg[22]  ( .D(\U16/Z_22 ), .CK(clock), .RN(n1531), 
        .Q(\U3/U1/DATA1_22 ), .QN(n34) );
  DFFR_X1 \scratchVal_FS_reg[22]  ( .D(\U20/Z_22 ), .CK(clock), .RN(n1532), 
        .Q(\U3/U1/DATA2_22 ) );
  DFFS_X2 \scratchVal_FS_reg[23]  ( .D(\U20/Z_23 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA2_23 ) );
  DFFR_X1 \scratchVal_Accum_reg[24]  ( .D(\U16/Z_24 ), .CK(clock), .RN(n1532), 
        .Q(\U3/U1/DATA1_24 ), .QN(n32) );
  DFFR_X1 \scratchVal_FS_reg[24]  ( .D(\U20/Z_24 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_24 ) );
  DFFS_X2 \scratchVal_FS_reg[25]  ( .D(\U20/Z_25 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA2_25 ) );
  DFFR_X1 \scratchVal_Accum_reg[26]  ( .D(\U16/Z_26 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA1_26 ), .QN(n30) );
  DFFR_X1 \scratchVal_FS_reg[26]  ( .D(\U20/Z_26 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA2_26 ) );
  DFFS_X2 \scratchVal_FS_reg[27]  ( .D(\U20/Z_27 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA2_27 ) );
  DFFR_X1 \scratchVal_Accum_reg[28]  ( .D(\U16/Z_28 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA1_28 ), .QN(n28) );
  DFFR_X1 \scratchVal_FS_reg[28]  ( .D(\U20/Z_28 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA2_28 ) );
  DFFS_X2 \scratchVal_FS_reg[29]  ( .D(\U20/Z_29 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA2_29 ) );
  DFFR_X1 \scratchVal_Accum_reg[30]  ( .D(\U16/Z_30 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA1_30 ), .QN(n26) );
  DFFR_X1 \scratchVal_FS_reg[30]  ( .D(\U20/Z_30 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_30 ) );
  DFFS_X2 \scratchVal_FS_reg[31]  ( .D(\U20/Z_31 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA2_31 ) );
  DFFR_X1 \scratchVal_FS_reg[32]  ( .D(\U20/Z_32 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_32 ) );
  DFFS_X2 \scratchVal_FS_reg[33]  ( .D(\U20/Z_33 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA2_33 ) );
  DFFR_X1 \scratchVal_Accum_reg[34]  ( .D(\U16/Z_34 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA1_34 ) );
  DFFR_X1 \scratchVal_FS_reg[34]  ( .D(\U20/Z_34 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_34 ) );
  DFFS_X2 \scratchVal_Accum_reg[35]  ( .D(\U16/Z_35 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA1_35 ), .QN(n21) );
  DFFR_X1 \scratchVal_FS_reg[9]  ( .D(\U20/Z_9 ), .CK(clock), .RN(n1535), .Q(
        \U3/U1/DATA2_9 ) );
  DFFR_X1 \scratchVal_FS_reg[8]  ( .D(\U20/Z_8 ), .CK(clock), .RN(n1534), .Q(
        \U3/U1/DATA2_8 ) );
  DFFR_X1 \scratchVal_FS_reg[7]  ( .D(\U20/Z_7 ), .CK(clock), .RN(n1535), .Q(
        \U3/U1/DATA2_7 ) );
  DFFR_X1 \scratchVal_FS_reg[6]  ( .D(\U20/Z_6 ), .CK(clock), .RN(n1534), .Q(
        \U3/U1/DATA2_6 ) );
  DFFR_X1 \scratchVal_FS_reg[5]  ( .D(\U20/Z_5 ), .CK(clock), .RN(n1535), .Q(
        \U3/U1/DATA2_5 ) );
  DFFR_X1 \scratchVal_FS_reg[4]  ( .D(\U20/Z_4 ), .CK(clock), .RN(n1534), .Q(
        \U3/U1/DATA2_4 ) );
  DFFR_X1 \scratchVal_FS_reg[3]  ( .D(\U20/Z_3 ), .CK(clock), .RN(n1534), .Q(
        \U3/U1/DATA2_3 ) );
  DFFR_X1 \scratchVal_FS_reg[2]  ( .D(\U20/Z_2 ), .CK(clock), .RN(n1534), .Q(
        \U3/U1/DATA2_2 ) );
  DFFR_X1 \scratchVal_FS_reg[19]  ( .D(\U20/Z_19 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA2_19 ) );
  DFFR_X1 \scratchVal_FS_reg[18]  ( .D(\U20/Z_18 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA2_18 ) );
  DFFR_X1 \scratchVal_FS_reg[17]  ( .D(\U20/Z_17 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_17 ) );
  DFFR_X1 \scratchVal_FS_reg[16]  ( .D(\U20/Z_16 ), .CK(clock), .RN(n1530), 
        .Q(\U3/U1/DATA2_16 ) );
  DFFR_X1 \scratchVal_FS_reg[15]  ( .D(\U20/Z_15 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_15 ) );
  DFFR_X1 \scratchVal_FS_reg[14]  ( .D(\U20/Z_14 ), .CK(clock), .RN(n1534), 
        .Q(\U3/U1/DATA2_14 ) );
  DFFR_X1 \scratchVal_FS_reg[13]  ( .D(\U20/Z_13 ), .CK(clock), .RN(rst_n), 
        .Q(\U3/U1/DATA2_13 ) );
  DFFR_X1 \scratchVal_FS_reg[12]  ( .D(\U20/Z_12 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_12 ) );
  DFFR_X1 \scratchVal_FS_reg[11]  ( .D(\U20/Z_11 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_11 ) );
  DFFR_X1 \scratchVal_FS_reg[10]  ( .D(\U20/Z_10 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA2_10 ) );
  DFFR_X1 \scratchVal_FS_reg[1]  ( .D(\U20/Z_1 ), .CK(clock), .RN(rst_n), .Q(
        \U3/U1/DATA2_1 ) );
  DFFS_X2 \scratchVal_FS_reg[35]  ( .D(\U20/Z_35 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA2_35 ) );
  AOI221_X2 U266 ( .B1(n1527), .B2(\U35/DATA2_34 ), .C1(n1454), .C2(
        \U35/DATA2_66 ), .A(n1836), .ZN(n239) );
  NAND2_X2 U268 ( .A1(n242), .A2(n243), .ZN(n219) );
  OAI22_X2 U271 ( .A1(n244), .A2(n121), .B1(\U15/DATA1_4 ), .B2(n245), .ZN(
        n220) );
  AOI221_X2 U272 ( .B1(\U35/DATA2_42 ), .B2(n1527), .C1(\U35/DATA1_10 ), .C2(
        n1454), .A(n1834), .ZN(n245) );
  AOI221_X2 U274 ( .B1(\U35/DATA2_58 ), .B2(n1527), .C1(\U35/DATA1_26 ), .C2(
        n1454), .A(n1833), .ZN(n244) );
  OAI22_X2 U277 ( .A1(n248), .A2(n121), .B1(\U15/DATA1_4 ), .B2(n249), .ZN(
        n190) );
  AOI221_X2 U278 ( .B1(\U35/DATA2_46 ), .B2(n1527), .C1(\U35/DATA1_14 ), .C2(
        n1454), .A(n1832), .ZN(n249) );
  AOI221_X2 U280 ( .B1(\U35/DATA2_62 ), .B2(n1527), .C1(\U35/DATA1_30 ), .C2(
        n1454), .A(n1831), .ZN(n248) );
  NAND2_X2 U282 ( .A1(n252), .A2(n253), .ZN(n191) );
  AOI221_X2 U285 ( .B1(\U35/DATA1_38 ), .B2(n1452), .C1(\U35/DATA2_6 ), .C2(
        n1451), .A(n1840), .ZN(n254) );
  AOI221_X2 U289 ( .B1(n1527), .B2(\U35/DATA2_32 ), .C1(n1454), .C2(
        \U35/DATA2_64 ), .A(n1829), .ZN(n257) );
  OAI22_X2 U293 ( .A1(n262), .A2(n121), .B1(\U15/DATA1_4 ), .B2(n263), .ZN(
        n261) );
  AOI221_X2 U294 ( .B1(\U35/DATA2_40 ), .B2(n1527), .C1(\U35/DATA1_8 ), .C2(
        n1454), .A(n1828), .ZN(n263) );
  AOI221_X2 U296 ( .B1(\U35/DATA2_56 ), .B2(n1527), .C1(\U35/DATA1_24 ), .C2(
        n1454), .A(n1827), .ZN(n262) );
  OAI22_X2 U299 ( .A1(n266), .A2(n121), .B1(\U15/DATA1_4 ), .B2(n267), .ZN(
        n205) );
  AOI221_X2 U300 ( .B1(\U35/DATA2_44 ), .B2(n1527), .C1(\U35/DATA1_12 ), .C2(
        n1454), .A(n1826), .ZN(n267) );
  AOI221_X2 U302 ( .B1(\U35/DATA2_60 ), .B2(n1527), .C1(\U35/DATA1_28 ), .C2(
        n1454), .A(n1825), .ZN(n266) );
  NAND2_X2 U304 ( .A1(n270), .A2(n271), .ZN(n207) );
  AOI221_X2 U307 ( .B1(\U35/DATA1_36 ), .B2(n1452), .C1(\U35/DATA2_4 ), .C2(
        n1451), .A(n1839), .ZN(n272) );
  OAI22_X2 U312 ( .A1(n278), .A2(n121), .B1(\U15/DATA1_4 ), .B2(n279), .ZN(
        n277) );
  AOI221_X2 U313 ( .B1(\U35/DATA2_45 ), .B2(n1527), .C1(\U35/DATA1_13 ), .C2(
        n1454), .A(n1823), .ZN(n279) );
  AOI221_X2 U315 ( .B1(\U35/DATA2_61 ), .B2(n1527), .C1(\U35/DATA1_29 ), .C2(
        n1454), .A(n1822), .ZN(n278) );
  AOI221_X2 U319 ( .B1(\U35/DATA1_37 ), .B2(n1452), .C1(\U35/DATA2_5 ), .C2(
        n1451), .A(n1838), .ZN(n276) );
  OAI22_X2 U322 ( .A1(n287), .A2(n121), .B1(\U15/DATA1_4 ), .B2(n288), .ZN(
        n286) );
  AOI221_X2 U323 ( .B1(\U35/DATA2_41 ), .B2(n1527), .C1(\U35/DATA1_9 ), .C2(
        n1454), .A(n1821), .ZN(n288) );
  AOI221_X2 U325 ( .B1(\U35/DATA2_57 ), .B2(n1527), .C1(\U35/DATA1_25 ), .C2(
        n1454), .A(n1820), .ZN(n287) );
  AOI221_X2 U329 ( .B1(\U35/DATA1_33 ), .B2(n1452), .C1(\U35/DATA2_1 ), .C2(
        n1451), .A(n1837), .ZN(n285) );
  AOI221_X2 U333 ( .B1(n1527), .B2(\U35/DATA2_35 ), .C1(n1454), .C2(
        \U35/DATA2_67 ), .A(n1819), .ZN(n295) );
  NOR2_X2 U335 ( .A1(\U15/DATA1_3 ), .A2(\U15/DATA1_4 ), .ZN(n238) );
  NAND2_X2 U336 ( .A1(n297), .A2(n298), .ZN(n214) );
  NOR2_X2 U339 ( .A1(n121), .A2(\U15/DATA1_3 ), .ZN(n237) );
  OAI22_X2 U340 ( .A1(n299), .A2(n121), .B1(\U15/DATA1_4 ), .B2(n300), .ZN(
        n213) );
  AOI221_X2 U341 ( .B1(\U35/DATA2_43 ), .B2(n1527), .C1(\U35/DATA1_11 ), .C2(
        n1454), .A(n1817), .ZN(n300) );
  AOI221_X2 U343 ( .B1(\U35/DATA2_59 ), .B2(n1527), .C1(\U35/DATA1_27 ), .C2(
        n1454), .A(n1816), .ZN(n299) );
  NOR2_X2 U361 ( .A1(n115), .A2(\U15/DATA1_6 ), .ZN(n192) );
  NAND4_X2 U422 ( .A1(n347), .A2(n348), .A3(n349), .A4(n350), .ZN(n346) );
  NOR4_X2 U423 ( .A1(\U28/DATA2_34 ), .A2(\U28/DATA2_32 ), .A3(\U28/DATA2_30 ), 
        .A4(\U28/DATA2_28 ), .ZN(n350) );
  NOR4_X2 U424 ( .A1(\U28/DATA2_26 ), .A2(\U28/DATA2_24 ), .A3(\U28/DATA2_22 ), 
        .A4(\U28/DATA2_20 ), .ZN(n349) );
  AND4_X2 U425 ( .A1(\U28/DATA2_27 ), .A2(\U28/DATA2_25 ), .A3(\U28/DATA2_23 ), 
        .A4(\U28/DATA2_21 ), .ZN(n348) );
  AND4_X2 U426 ( .A1(\U28/DATA2_35 ), .A2(\U28/DATA2_33 ), .A3(\U28/DATA2_31 ), 
        .A4(\U28/DATA2_29 ), .ZN(n347) );
  NOR4_X2 U428 ( .A1(input_done), .A2(n355), .A3(n356), .A4(n357), .ZN(n354)
         );
  NOR4_X2 U432 ( .A1(n358), .A2(n359), .A3(n360), .A4(n361), .ZN(n353) );
  NOR4_X2 U447 ( .A1(n370), .A2(n371), .A3(n372), .A4(n373), .ZN(n344) );
  NAND4_X2 U448 ( .A1(\U28/DATA1_35 ), .A2(\U28/DATA1_33 ), .A3(\U28/DATA1_31 ), .A4(\U28/DATA1_29 ), .ZN(n373) );
  NAND2_X2 U496 ( .A1(n1460), .A2(n147), .ZN(\U14/Z_0 ) );
  NOR2_X2 U506 ( .A1(n121), .A2(n123), .ZN(n208) );
  AND2_X1 U572 ( .A1(\U26/DATA1_0 ), .A2(n1521), .ZN(\U26/Z_0 ) );
  AND2_X1 U573 ( .A1(\U25/DATA1_0 ), .A2(n1521), .ZN(\U25/Z_0 ) );
  AND2_X1 U574 ( .A1(n259), .A2(n260), .ZN(n233) );
  AND2_X1 U575 ( .A1(n282), .A2(n283), .ZN(n201) );
  AND2_X1 U576 ( .A1(n291), .A2(n292), .ZN(n227) );
  AND2_X1 U577 ( .A1(n303), .A2(n304), .ZN(n212) );
  AND2_X1 U578 ( .A1(\U23/DATA1_0 ), .A2(n1521), .ZN(\U23/Z_0 ) );
  AND2_X1 U579 ( .A1(\U22/DATA1_0 ), .A2(n1521), .ZN(\U22/Z_0 ) );
  OR4_X1 U590 ( .A1(\U28/DATA1_30 ), .A2(\U28/DATA1_28 ), .A3(\U28/DATA1_34 ), 
        .A4(\U28/DATA1_32 ), .ZN(n370) );
  AND2_X1 U591 ( .A1(\U19/DATA1_0 ), .A2(n1521), .ZN(\U19/Z_0 ) );
  DFFR_X2 \pipelineCounter_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n1529), .Q(
        \U15/DATA1_3 ), .QN(n123) );
  DFFR_X2 \pipelineCounter_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(n1529), .Q(
        \U15/DATA1_4 ), .QN(n121) );
  DFFS_X2 \scratchVal_Accum_reg[33]  ( .D(n1514), .CK(clock), .SN(rst_n), .Q(
        \U3/U1/DATA1_33 ), .QN(n23) );
  DFFR_X2 \readInitial_Accum_reg[5]  ( .D(\U17/Z_5 ), .CK(clock), .RN(n1531), 
        .Q(\eq_122/B[5] ), .QN(n1509) );
  DFFR_X2 \readInitial_FS_reg[6]  ( .D(\U21/Z_6 ), .CK(clock), .RN(n1531), .Q(
        \U17/DATA1_6 ), .QN(n1540) );
  DFFR_X2 \scratchVal_Accum_reg[32]  ( .D(\U16/Z_32 ), .CK(clock), .RN(n1535), 
        .Q(\U3/U1/DATA1_32 ), .QN(n24) );
  DFFR_X1 \scratchVal_Accum_reg[16]  ( .D(\U16/Z_16 ), .CK(clock), .RN(n1533), 
        .Q(\U3/U1/DATA1_16 ), .QN(n40) );
  DFFR_X2 \memoryCounter_reg[0]  ( .D(n421), .CK(clock), .RN(n1533), .Q(
        \U5/DATA1_0 ), .QN(n128) );
  DFFR_X2 \memoryCounter_reg[15]  ( .D(n420), .CK(clock), .RN(n1531), .Q(
        \U5/DATA1_15 ), .QN(n127) );
  DFFR_X2 \readInitial_FS_reg[4]  ( .D(\U21/Z_4 ), .CK(clock), .RN(n1531), 
        .QN(n1481) );
  DFFR_X2 \readInitial_Accum_reg[1]  ( .D(\U17/Z_1 ), .CK(clock), .RN(n1532), 
        .Q(\eq_122/B[1] ), .QN(n1479) );
  DFFR_X2 \readInitial_Accum_reg[0]  ( .D(\U17/Z_0 ), .CK(clock), .RN(n1532), 
        .Q(\eq_122/B[0] ), .QN(n1477) );
  DFF_X2 \m3WriteAddr_reg[14]  ( .D(\U5/DATA1_14 ), .CK(clock), .Q(
        m3WriteAddr[14]) );
  DFF_X2 \m3WriteAddr_reg[13]  ( .D(\U5/DATA1_13 ), .CK(clock), .Q(
        m3WriteAddr[13]) );
  DFF_X2 \m3WriteAddr_reg[12]  ( .D(\U5/DATA1_12 ), .CK(clock), .Q(
        m3WriteAddr[12]) );
  DFF_X2 \m3WriteAddr_reg[11]  ( .D(\U5/DATA1_11 ), .CK(clock), .Q(
        m3WriteAddr[11]) );
  DFF_X2 \m3WriteAddr_reg[10]  ( .D(\U5/DATA1_10 ), .CK(clock), .Q(
        m3WriteAddr[10]) );
  DFF_X2 \m3WriteAddr_reg[9]  ( .D(\U5/DATA1_9 ), .CK(clock), .Q(
        m3WriteAddr[9]) );
  DFF_X2 \m3WriteAddr_reg[8]  ( .D(\U5/DATA1_8 ), .CK(clock), .Q(
        m3WriteAddr[8]) );
  DFF_X2 \m3WriteAddr_reg[7]  ( .D(\U5/DATA1_7 ), .CK(clock), .Q(
        m3WriteAddr[7]) );
  DFF_X2 \m3WriteAddr_reg[6]  ( .D(\U5/DATA1_6 ), .CK(clock), .Q(
        m3WriteAddr[6]) );
  DFF_X2 \m3WriteAddr_reg[5]  ( .D(\U5/DATA1_5 ), .CK(clock), .Q(
        m3WriteAddr[5]) );
  DFF_X2 \m3WriteAddr_reg[4]  ( .D(\U5/DATA1_4 ), .CK(clock), .Q(
        m3WriteAddr[4]) );
  DFF_X2 \m3WriteAddr_reg[3]  ( .D(\U5/DATA1_3 ), .CK(clock), .Q(
        m3WriteAddr[3]) );
  DFF_X2 \m3WriteAddr_reg[2]  ( .D(\U5/DATA1_2 ), .CK(clock), .Q(
        m3WriteAddr[2]) );
  DFF_X2 \m3WriteAddr_reg[1]  ( .D(\U5/DATA1_1 ), .CK(clock), .Q(
        m3WriteAddr[1]) );
  DFF_X2 m3WE_reg ( .D(\U22/DATA1_0 ), .CK(clock), .Q(m3WE) );
  DFF_X2 \m3WriteAddr_reg[0]  ( .D(\U5/DATA1_0 ), .CK(clock), .Q(
        m3WriteAddr[0]) );
  DFF_X2 \m3WriteBus_reg[0]  ( .D(\U35/DATA2_0 ), .CK(clock), .Q(m3WriteBus[0]) );
  DFF_X2 \m3WriteBus_reg[1]  ( .D(\U35/DATA2_1 ), .CK(clock), .Q(m3WriteBus[1]) );
  DFF_X2 \m3WriteBus_reg[2]  ( .D(\U35/DATA2_2 ), .CK(clock), .Q(m3WriteBus[2]) );
  DFF_X2 \m3WriteBus_reg[3]  ( .D(\U35/DATA2_3 ), .CK(clock), .Q(m3WriteBus[3]) );
  DFF_X2 \m3WriteBus_reg[4]  ( .D(\U35/DATA2_4 ), .CK(clock), .Q(m3WriteBus[4]) );
  DFF_X2 \m3WriteBus_reg[5]  ( .D(\U35/DATA2_5 ), .CK(clock), .Q(m3WriteBus[5]) );
  DFF_X2 \m3WriteBus_reg[6]  ( .D(\U35/DATA2_6 ), .CK(clock), .Q(m3WriteBus[6]) );
  DFF_X2 \m3WriteBus_reg[7]  ( .D(\U35/DATA2_7 ), .CK(clock), .Q(m3WriteBus[7]) );
  DFF_X2 \m3WriteBus_reg[8]  ( .D(\U35/DATA2_8 ), .CK(clock), .Q(m3WriteBus[8]) );
  DFF_X2 \m3WriteBus_reg[9]  ( .D(\U35/DATA2_9 ), .CK(clock), .Q(m3WriteBus[9]) );
  DFF_X2 \m3WriteBus_reg[10]  ( .D(\U35/DATA2_10 ), .CK(clock), .Q(
        m3WriteBus[10]) );
  DFF_X2 \m3WriteBus_reg[11]  ( .D(\U35/DATA2_11 ), .CK(clock), .Q(
        m3WriteBus[11]) );
  DFF_X2 \m3WriteBus_reg[12]  ( .D(\U35/DATA2_12 ), .CK(clock), .Q(
        m3WriteBus[12]) );
  DFF_X2 \m3WriteBus_reg[13]  ( .D(\U35/DATA2_13 ), .CK(clock), .Q(
        m3WriteBus[13]) );
  DFF_X2 \m3WriteBus_reg[14]  ( .D(\U35/DATA2_14 ), .CK(clock), .Q(
        m3WriteBus[14]) );
  DFF_X2 \m3WriteBus_reg[15]  ( .D(\U35/DATA2_15 ), .CK(clock), .Q(
        m3WriteBus[15]) );
  DFF_X2 \m3WriteBus_reg[16]  ( .D(\U35/DATA2_16 ), .CK(clock), .Q(
        m3WriteBus[16]) );
  DFF_X2 \m3WriteBus_reg[17]  ( .D(\U35/DATA2_17 ), .CK(clock), .Q(
        m3WriteBus[17]) );
  DFF_X2 \m3WriteBus_reg[18]  ( .D(\U35/DATA2_18 ), .CK(clock), .Q(
        m3WriteBus[18]) );
  DFF_X2 \m3WriteBus_reg[19]  ( .D(\U35/DATA2_19 ), .CK(clock), .Q(
        m3WriteBus[19]) );
  DFF_X2 \m3WriteBus_reg[20]  ( .D(\U35/DATA2_20 ), .CK(clock), .Q(
        m3WriteBus[20]) );
  DFF_X2 \m3WriteBus_reg[21]  ( .D(\U35/DATA2_21 ), .CK(clock), .Q(
        m3WriteBus[21]) );
  DFF_X2 \m3WriteBus_reg[22]  ( .D(\U35/DATA2_22 ), .CK(clock), .Q(
        m3WriteBus[22]) );
  DFF_X2 \m3WriteBus_reg[23]  ( .D(\U35/DATA2_23 ), .CK(clock), .Q(
        m3WriteBus[23]) );
  DFF_X2 \m3WriteBus_reg[24]  ( .D(\U35/DATA2_24 ), .CK(clock), .Q(
        m3WriteBus[24]) );
  DFF_X2 \m3WriteBus_reg[25]  ( .D(\U35/DATA2_25 ), .CK(clock), .Q(
        m3WriteBus[25]) );
  DFF_X2 \m3WriteBus_reg[26]  ( .D(\U35/DATA2_26 ), .CK(clock), .Q(
        m3WriteBus[26]) );
  DFF_X2 \m3WriteBus_reg[27]  ( .D(\U35/DATA2_27 ), .CK(clock), .Q(
        m3WriteBus[27]) );
  DFF_X2 \m3WriteBus_reg[28]  ( .D(\U35/DATA2_28 ), .CK(clock), .Q(
        m3WriteBus[28]) );
  DFF_X2 \m3WriteBus_reg[29]  ( .D(\U35/DATA2_29 ), .CK(clock), .Q(
        m3WriteBus[29]) );
  DFF_X2 \m3WriteBus_reg[30]  ( .D(\U35/DATA2_30 ), .CK(clock), .Q(
        m3WriteBus[30]) );
  DFF_X2 \m3WriteBus_reg[31]  ( .D(\U35/DATA2_31 ), .CK(clock), .Q(
        m3WriteBus[31]) );
  DFF_X2 \m3WriteBus_reg[32]  ( .D(\U35/DATA2_32 ), .CK(clock), .Q(
        m3WriteBus[32]) );
  DFF_X2 \m3WriteBus_reg[33]  ( .D(\U35/DATA2_33 ), .CK(clock), .Q(
        m3WriteBus[33]) );
  DFF_X2 \m3WriteBus_reg[34]  ( .D(\U35/DATA2_34 ), .CK(clock), .Q(
        m3WriteBus[34]) );
  DFF_X2 \m3WriteBus_reg[35]  ( .D(\U35/DATA2_35 ), .CK(clock), .Q(
        m3WriteBus[35]) );
  DFF_X2 \m3WriteBus_reg[36]  ( .D(\U35/DATA2_36 ), .CK(clock), .Q(
        m3WriteBus[36]) );
  DFF_X2 \m3WriteBus_reg[37]  ( .D(\U35/DATA2_37 ), .CK(clock), .Q(
        m3WriteBus[37]) );
  DFF_X2 \m3WriteBus_reg[38]  ( .D(\U35/DATA2_38 ), .CK(clock), .Q(
        m3WriteBus[38]) );
  DFF_X2 \m3WriteBus_reg[39]  ( .D(\U35/DATA2_39 ), .CK(clock), .Q(
        m3WriteBus[39]) );
  DFF_X2 \m3WriteBus_reg[40]  ( .D(\U35/DATA2_40 ), .CK(clock), .Q(
        m3WriteBus[40]) );
  DFF_X2 \m3WriteBus_reg[41]  ( .D(\U35/DATA2_41 ), .CK(clock), .Q(
        m3WriteBus[41]) );
  DFF_X2 \m3WriteBus_reg[42]  ( .D(\U35/DATA2_42 ), .CK(clock), .Q(
        m3WriteBus[42]) );
  DFF_X2 \m3WriteBus_reg[43]  ( .D(\U35/DATA2_43 ), .CK(clock), .Q(
        m3WriteBus[43]) );
  DFF_X2 \m3WriteBus_reg[44]  ( .D(\U35/DATA2_44 ), .CK(clock), .Q(
        m3WriteBus[44]) );
  DFF_X2 \m3WriteBus_reg[45]  ( .D(\U35/DATA2_45 ), .CK(clock), .Q(
        m3WriteBus[45]) );
  DFF_X2 \m3WriteBus_reg[46]  ( .D(\U35/DATA2_46 ), .CK(clock), .Q(
        m3WriteBus[46]) );
  DFF_X2 \m3WriteBus_reg[47]  ( .D(\U35/DATA2_47 ), .CK(clock), .Q(
        m3WriteBus[47]) );
  DFF_X2 \m3WriteBus_reg[48]  ( .D(\U35/DATA2_48 ), .CK(clock), .Q(
        m3WriteBus[48]) );
  DFF_X2 \m3WriteBus_reg[49]  ( .D(\U35/DATA2_49 ), .CK(clock), .Q(
        m3WriteBus[49]) );
  DFF_X2 \m3WriteBus_reg[50]  ( .D(\U35/DATA2_50 ), .CK(clock), .Q(
        m3WriteBus[50]) );
  DFF_X2 \m3WriteBus_reg[51]  ( .D(\U35/DATA2_51 ), .CK(clock), .Q(
        m3WriteBus[51]) );
  DFF_X2 \m3WriteBus_reg[52]  ( .D(\U35/DATA2_52 ), .CK(clock), .Q(
        m3WriteBus[52]) );
  DFF_X2 \m3WriteBus_reg[53]  ( .D(\U35/DATA2_53 ), .CK(clock), .Q(
        m3WriteBus[53]) );
  DFF_X2 \m3WriteBus_reg[54]  ( .D(\U35/DATA2_54 ), .CK(clock), .Q(
        m3WriteBus[54]) );
  DFF_X2 \m3WriteBus_reg[55]  ( .D(\U35/DATA2_55 ), .CK(clock), .Q(
        m3WriteBus[55]) );
  DFF_X2 \m3WriteBus_reg[56]  ( .D(\U35/DATA2_56 ), .CK(clock), .Q(
        m3WriteBus[56]) );
  DFF_X2 \m3WriteBus_reg[57]  ( .D(\U35/DATA2_57 ), .CK(clock), .Q(
        m3WriteBus[57]) );
  DFF_X2 \m3WriteBus_reg[58]  ( .D(\U35/DATA2_58 ), .CK(clock), .Q(
        m3WriteBus[58]) );
  DFF_X2 \m3WriteBus_reg[59]  ( .D(\U35/DATA2_59 ), .CK(clock), .Q(
        m3WriteBus[59]) );
  DFF_X2 \m3WriteBus_reg[60]  ( .D(\U35/DATA2_60 ), .CK(clock), .Q(
        m3WriteBus[60]) );
  DFF_X2 \m3WriteBus_reg[61]  ( .D(\U35/DATA2_61 ), .CK(clock), .Q(
        m3WriteBus[61]) );
  DFF_X2 \m3WriteBus_reg[62]  ( .D(\U35/DATA2_62 ), .CK(clock), .Q(
        m3WriteBus[62]) );
  DFF_X2 \m3WriteBus_reg[63]  ( .D(\U35/DATA2_63 ), .CK(clock), .Q(
        m3WriteBus[63]) );
  DFF_X2 \m3WriteBus_reg[64]  ( .D(\U35/DATA2_64 ), .CK(clock), .Q(
        m3WriteBus[64]) );
  DFF_X2 \m3WriteBus_reg[65]  ( .D(\U35/DATA2_65 ), .CK(clock), .Q(
        m3WriteBus[65]) );
  DFF_X2 \m3WriteBus_reg[66]  ( .D(\U35/DATA2_66 ), .CK(clock), .Q(
        m3WriteBus[66]) );
  DFF_X2 \m3WriteBus_reg[67]  ( .D(\U35/DATA2_67 ), .CK(clock), .Q(
        m3WriteBus[67]) );
  DFF_X2 \m3WriteBus_reg[68]  ( .D(\U35/DATA2_68 ), .CK(clock), .Q(
        m3WriteBus[68]) );
  DFF_X2 \m3WriteBus_reg[69]  ( .D(\U35/DATA2_69 ), .CK(clock), .Q(
        m3WriteBus[69]) );
  DFF_X2 \m3WriteBus_reg[70]  ( .D(\U35/DATA2_70 ), .CK(clock), .Q(
        m3WriteBus[70]) );
  DFF_X2 \m3WriteBus_reg[71]  ( .D(\U35/DATA1_7 ), .CK(clock), .Q(
        m3WriteBus[71]) );
  DFF_X2 \m3WriteBus_reg[72]  ( .D(\U35/DATA1_8 ), .CK(clock), .Q(
        m3WriteBus[72]) );
  DFF_X2 \m3WriteBus_reg[73]  ( .D(\U35/DATA1_9 ), .CK(clock), .Q(
        m3WriteBus[73]) );
  DFF_X2 \m3WriteBus_reg[74]  ( .D(\U35/DATA1_10 ), .CK(clock), .Q(
        m3WriteBus[74]) );
  DFF_X2 \m3WriteBus_reg[75]  ( .D(\U35/DATA1_11 ), .CK(clock), .Q(
        m3WriteBus[75]) );
  DFF_X2 \m3WriteBus_reg[76]  ( .D(\U35/DATA1_12 ), .CK(clock), .Q(
        m3WriteBus[76]) );
  DFF_X2 \m3WriteBus_reg[77]  ( .D(\U35/DATA1_13 ), .CK(clock), .Q(
        m3WriteBus[77]) );
  DFF_X2 \m3WriteBus_reg[78]  ( .D(\U35/DATA1_14 ), .CK(clock), .Q(
        m3WriteBus[78]) );
  DFF_X2 \m3WriteBus_reg[79]  ( .D(\U35/DATA1_15 ), .CK(clock), .Q(
        m3WriteBus[79]) );
  DFF_X2 \m3WriteBus_reg[80]  ( .D(\U35/DATA1_16 ), .CK(clock), .Q(
        m3WriteBus[80]) );
  DFF_X2 \m3WriteBus_reg[81]  ( .D(\U35/DATA1_17 ), .CK(clock), .Q(
        m3WriteBus[81]) );
  DFF_X2 \m3WriteBus_reg[82]  ( .D(\U35/DATA1_18 ), .CK(clock), .Q(
        m3WriteBus[82]) );
  DFF_X2 \m3WriteBus_reg[83]  ( .D(\U35/DATA1_19 ), .CK(clock), .Q(
        m3WriteBus[83]) );
  DFF_X2 \m3WriteBus_reg[84]  ( .D(\U35/DATA1_20 ), .CK(clock), .Q(
        m3WriteBus[84]) );
  DFF_X2 \m3WriteBus_reg[85]  ( .D(\U35/DATA1_21 ), .CK(clock), .Q(
        m3WriteBus[85]) );
  DFF_X2 \m3WriteBus_reg[86]  ( .D(\U35/DATA1_22 ), .CK(clock), .Q(
        m3WriteBus[86]) );
  DFF_X2 \m3WriteBus_reg[87]  ( .D(\U35/DATA1_23 ), .CK(clock), .Q(
        m3WriteBus[87]) );
  DFF_X2 \m3WriteBus_reg[88]  ( .D(\U35/DATA1_24 ), .CK(clock), .Q(
        m3WriteBus[88]) );
  DFF_X2 \m3WriteBus_reg[89]  ( .D(\U35/DATA1_25 ), .CK(clock), .Q(
        m3WriteBus[89]) );
  DFF_X2 \m3WriteBus_reg[90]  ( .D(\U35/DATA1_26 ), .CK(clock), .Q(
        m3WriteBus[90]) );
  DFF_X2 \m3WriteBus_reg[91]  ( .D(\U35/DATA1_27 ), .CK(clock), .Q(
        m3WriteBus[91]) );
  DFF_X2 \m3WriteBus_reg[92]  ( .D(\U35/DATA1_28 ), .CK(clock), .Q(
        m3WriteBus[92]) );
  DFF_X2 \m3WriteBus_reg[93]  ( .D(\U35/DATA1_29 ), .CK(clock), .Q(
        m3WriteBus[93]) );
  DFF_X2 \m3WriteBus_reg[94]  ( .D(\U35/DATA1_30 ), .CK(clock), .Q(
        m3WriteBus[94]) );
  DFF_X2 \m3WriteBus_reg[95]  ( .D(\U35/DATA1_31 ), .CK(clock), .Q(
        m3WriteBus[95]) );
  DFF_X2 \m3WriteBus_reg[96]  ( .D(\U35/DATA1_32 ), .CK(clock), .Q(
        m3WriteBus[96]) );
  DFF_X2 \m3WriteBus_reg[97]  ( .D(\U35/DATA1_33 ), .CK(clock), .Q(
        m3WriteBus[97]) );
  DFF_X2 \m3WriteBus_reg[98]  ( .D(\U35/DATA1_34 ), .CK(clock), .Q(
        m3WriteBus[98]) );
  DFF_X2 \m3WriteBus_reg[99]  ( .D(\U35/DATA1_35 ), .CK(clock), .Q(
        m3WriteBus[99]) );
  DFF_X2 \m3WriteBus_reg[100]  ( .D(\U35/DATA1_36 ), .CK(clock), .Q(
        m3WriteBus[100]) );
  DFF_X2 \m3WriteBus_reg[101]  ( .D(\U35/DATA1_37 ), .CK(clock), .Q(
        m3WriteBus[101]) );
  DFF_X2 \m3WriteBus_reg[102]  ( .D(\U35/DATA1_38 ), .CK(clock), .Q(
        m3WriteBus[102]) );
  DFF_X2 \m3WriteBus_reg[103]  ( .D(\U35/DATA1_39 ), .CK(clock), .Q(
        m3WriteBus[103]) );
  DFF_X2 \m3WriteBus_reg[104]  ( .D(\U35/DATA1_40 ), .CK(clock), .Q(
        m3WriteBus[104]) );
  DFF_X2 \m3WriteBus_reg[105]  ( .D(\U35/DATA1_41 ), .CK(clock), .Q(
        m3WriteBus[105]) );
  DFF_X2 \m3WriteBus_reg[106]  ( .D(\U35/DATA1_42 ), .CK(clock), .Q(
        m3WriteBus[106]) );
  DFF_X2 \m3WriteBus_reg[107]  ( .D(\U35/DATA1_43 ), .CK(clock), .Q(
        m3WriteBus[107]) );
  DFF_X2 \m3WriteBus_reg[108]  ( .D(\U35/DATA1_44 ), .CK(clock), .Q(
        m3WriteBus[108]) );
  DFF_X2 \m3WriteBus_reg[109]  ( .D(\U35/DATA1_45 ), .CK(clock), .Q(
        m3WriteBus[109]) );
  DFF_X2 \m3WriteBus_reg[110]  ( .D(\U35/DATA1_46 ), .CK(clock), .Q(
        m3WriteBus[110]) );
  DFF_X2 \m3WriteBus_reg[111]  ( .D(\U35/DATA1_47 ), .CK(clock), .Q(
        m3WriteBus[111]) );
  DFF_X2 \m3WriteBus_reg[112]  ( .D(\U35/DATA1_48 ), .CK(clock), .Q(
        m3WriteBus[112]) );
  DFF_X2 \m3WriteBus_reg[113]  ( .D(\U35/DATA1_49 ), .CK(clock), .Q(
        m3WriteBus[113]) );
  DFF_X2 \m3WriteBus_reg[114]  ( .D(\U35/DATA1_50 ), .CK(clock), .Q(
        m3WriteBus[114]) );
  DFF_X2 \m3WriteBus_reg[115]  ( .D(\U35/DATA1_51 ), .CK(clock), .Q(
        m3WriteBus[115]) );
  DFF_X2 \m3WriteBus_reg[116]  ( .D(\U35/DATA1_52 ), .CK(clock), .Q(
        m3WriteBus[116]) );
  DFF_X2 \m3WriteBus_reg[117]  ( .D(\U35/DATA1_53 ), .CK(clock), .Q(
        m3WriteBus[117]) );
  DFF_X2 \m3WriteBus_reg[118]  ( .D(\U35/DATA1_54 ), .CK(clock), .Q(
        m3WriteBus[118]) );
  DFF_X2 \m3WriteBus_reg[119]  ( .D(\U35/DATA1_55 ), .CK(clock), .Q(
        m3WriteBus[119]) );
  DFF_X2 \m3WriteBus_reg[120]  ( .D(\U35/DATA1_56 ), .CK(clock), .Q(
        m3WriteBus[120]) );
  DFF_X2 \m3WriteBus_reg[121]  ( .D(\U35/DATA1_57 ), .CK(clock), .Q(
        m3WriteBus[121]) );
  DFF_X2 \m3WriteBus_reg[122]  ( .D(\U35/DATA1_58 ), .CK(clock), .Q(
        m3WriteBus[122]) );
  DFF_X2 \m3WriteBus_reg[123]  ( .D(\U35/DATA1_59 ), .CK(clock), .Q(
        m3WriteBus[123]) );
  DFF_X2 \m3WriteBus_reg[124]  ( .D(\U35/DATA1_60 ), .CK(clock), .Q(
        m3WriteBus[124]) );
  DFF_X2 \m3WriteBus_reg[125]  ( .D(\U35/DATA1_61 ), .CK(clock), .Q(
        m3WriteBus[125]) );
  DFF_X2 \m3WriteBus_reg[126]  ( .D(\U35/DATA1_62 ), .CK(clock), .Q(
        m3WriteBus[126]) );
  DFF_X2 \m3WriteBus_reg[127]  ( .D(\U35/DATA1_63 ), .CK(clock), .Q(
        m3WriteBus[127]) );
  DFF_X2 \m3WriteAddr_reg[15]  ( .D(inputBaseOffset), .CK(clock), .Q(
        m3WriteAddr[15]) );
  DFFR_X1 \readInitial_FS_reg[3]  ( .D(\U21/Z_3 ), .CK(clock), .RN(n1531), .Q(
        n1450), .QN(n1474) );
  DFFR_X2 \scratchVal_Accum_reg[0]  ( .D(n1471), .CK(clock), .RN(rst_n), .Q(
        \U3/U1/DATA1_0 ), .QN(n57) );
  SDFFR_X1 \readInitial_FI_reg[7]  ( .D(start), .SI(1'b0), .SE(n212), .CK(
        clock), .RN(rst_n), .Q(\U21/DATA1_7 ), .QN(n1537) );
  DFFS_X2 \scratchVal_Accum_reg[29]  ( .D(n1469), .CK(clock), .SN(rst_n), .Q(
        \U3/U1/DATA1_29 ), .QN(n27) );
  DFFS_X2 \scratchVal_Accum_reg[23]  ( .D(n1468), .CK(clock), .SN(rst_n), .Q(
        \U3/U1/DATA1_23 ), .QN(n33) );
  DFFS_X2 \scratchVal_Accum_reg[25]  ( .D(n1467), .CK(clock), .SN(rst_n), .Q(
        \U3/U1/DATA1_25 ), .QN(n31) );
  DFFS_X2 \scratchVal_Accum_reg[27]  ( .D(n1466), .CK(clock), .SN(rst_n), .Q(
        \U3/U1/DATA1_27 ), .QN(n29) );
  DFFS_X2 \scratchVal_Accum_reg[21]  ( .D(n1465), .CK(clock), .SN(rst_n), .Q(
        \U3/U1/DATA1_21 ), .QN(n35) );
  DFFS_X2 \scratchVal_Accum_reg[31]  ( .D(n1464), .CK(clock), .SN(rst_n), .Q(
        \U3/U1/DATA1_31 ), .QN(n25) );
  DFF_X2 \m2WriteBus_reg[29]  ( .D(\U3/U1/DATA1_29 ), .CK(clock), .Q(
        \U28/DATA1_29 ) );
  DFF_X2 \m2WriteBus_reg[31]  ( .D(\U3/U1/DATA1_31 ), .CK(clock), .Q(
        \U28/DATA1_31 ) );
  DFF_X2 \m2WriteBus_reg[27]  ( .D(\U3/U1/DATA1_27 ), .CK(clock), .Q(
        \U28/DATA1_27 ) );
  DFF_X2 \m2WriteBus_reg[25]  ( .D(\U3/U1/DATA1_25 ), .CK(clock), .Q(
        \U28/DATA1_25 ) );
  DFF_X2 \m2WriteBus_reg[23]  ( .D(\U3/U1/DATA1_23 ), .CK(clock), .Q(
        \U28/DATA1_23 ) );
  DFF_X2 \m2WriteBus_reg[21]  ( .D(\U3/U1/DATA1_21 ), .CK(clock), .Q(
        \U28/DATA1_21 ) );
  DFF_X2 \m2WriteBus_reg[0]  ( .D(\U3/U1/DATA1_0 ), .CK(clock), .Q(
        \U28/DATA1_0 ), .QN(n1558) );
  DFF_X2 \m2WriteBus_reg[30]  ( .D(\U3/U1/DATA1_30 ), .CK(clock), .Q(
        \U28/DATA1_30 ) );
  DFF_X2 \m2WriteBus_reg[28]  ( .D(\U3/U1/DATA1_28 ), .CK(clock), .Q(
        \U28/DATA1_28 ) );
  DFF_X2 \m2WriteBus_reg[26]  ( .D(\U3/U1/DATA1_26 ), .CK(clock), .Q(
        \U28/DATA1_26 ), .QN(n1788) );
  DFF_X2 \m2WriteBus_reg[24]  ( .D(\U3/U1/DATA1_24 ), .CK(clock), .Q(
        \U28/DATA1_24 ), .QN(n1789) );
  DFF_X2 \m2WriteBus_reg[22]  ( .D(\U3/U1/DATA1_22 ), .CK(clock), .Q(
        \U28/DATA1_22 ), .QN(n1790) );
  DFF_X2 \m2WriteBus_reg[20]  ( .D(\U3/U1/DATA1_20 ), .CK(clock), .Q(
        \U28/DATA1_20 ), .QN(n1791) );
  DFF_X2 \m2WriteBus_reg[19]  ( .D(\U3/U1/DATA1_19 ), .CK(clock), .Q(
        \U28/DATA1_19 ), .QN(n1665) );
  DFF_X2 \m2WriteBus_reg[18]  ( .D(\U3/U1/DATA1_18 ), .CK(clock), .Q(
        \U28/DATA1_18 ), .QN(n1659) );
  DFF_X2 \m2WriteBus_reg[17]  ( .D(\U3/U1/DATA1_17 ), .CK(clock), .Q(
        \U28/DATA1_17 ), .QN(n1643) );
  DFF_X2 \m2WriteBus_reg[16]  ( .D(\U3/U1/DATA1_16 ), .CK(clock), .Q(
        \U28/DATA1_16 ), .QN(n1637) );
  DFF_X2 \m2WriteBus_reg[15]  ( .D(\U3/U1/DATA1_15 ), .CK(clock), .Q(
        \U28/DATA1_15 ), .QN(n1632) );
  DFF_X2 \m2WriteBus_reg[14]  ( .D(\U3/U1/DATA1_14 ), .CK(clock), .Q(
        \U28/DATA1_14 ), .QN(n1628) );
  DFF_X2 \m2WriteBus_reg[13]  ( .D(\U3/U1/DATA1_13 ), .CK(clock), .Q(
        \U28/DATA1_13 ), .QN(n1624) );
  DFF_X2 \m2WriteBus_reg[12]  ( .D(\U3/U1/DATA1_12 ), .CK(clock), .Q(
        \U28/DATA1_12 ), .QN(n1620) );
  DFF_X2 \m2WriteBus_reg[11]  ( .D(\U3/U1/DATA1_11 ), .CK(clock), .Q(
        \U28/DATA1_11 ), .QN(n1616) );
  DFF_X2 \m2WriteBus_reg[10]  ( .D(\U3/U1/DATA1_10 ), .CK(clock), .Q(
        \U28/DATA1_10 ), .QN(n1613) );
  DFF_X2 \m2WriteBus_reg[9]  ( .D(\U3/U1/DATA1_9 ), .CK(clock), .Q(
        \U28/DATA1_9 ), .QN(n1598) );
  DFF_X2 \m2WriteBus_reg[8]  ( .D(\U3/U1/DATA1_8 ), .CK(clock), .Q(
        \U28/DATA1_8 ), .QN(n1592) );
  DFF_X2 \m2WriteBus_reg[7]  ( .D(\U3/U1/DATA1_7 ), .CK(clock), .Q(
        \U28/DATA1_7 ), .QN(n1589) );
  DFF_X2 \m2WriteBus_reg[6]  ( .D(\U3/U1/DATA1_6 ), .CK(clock), .Q(
        \U28/DATA1_6 ), .QN(n1586) );
  DFF_X2 \m2WriteBus_reg[5]  ( .D(\U3/U1/DATA1_5 ), .CK(clock), .Q(
        \U28/DATA1_5 ), .QN(n1583) );
  DFF_X2 \m2WriteBus_reg[4]  ( .D(\U3/U1/DATA1_4 ), .CK(clock), .Q(
        \U28/DATA1_4 ), .QN(n1580) );
  DFF_X2 \m2WriteBus_reg[3]  ( .D(\U3/U1/DATA1_3 ), .CK(clock), .Q(
        \U28/DATA1_3 ), .QN(n1577) );
  DFF_X2 \m2WriteBus_reg[2]  ( .D(\U3/U1/DATA1_2 ), .CK(clock), .Q(
        \U28/DATA1_2 ), .QN(n1574) );
  DFF_X2 \m2WriteBus_reg[1]  ( .D(\U3/U1/DATA1_1 ), .CK(clock), .Q(
        \U28/DATA1_1 ), .QN(n1571) );
  DFF_X2 m2WE_reg ( .D(n501), .CK(clock), .Q(m2WE) );
  DFF_X2 input_done_reg ( .D(n448), .CK(clock), .Q(input_done) );
  DFF_X2 \m2WriteBus_reg[32]  ( .D(\U3/U1/DATA1_32 ), .CK(clock), .Q(
        \U28/DATA1_32 ) );
  DFF_X2 \m2WriteBus_reg[34]  ( .D(\U3/U1/DATA1_34 ), .CK(clock), .Q(
        \U28/DATA1_34 ) );
  DFF_X2 \m2WriteBus_reg[35]  ( .D(\U3/U1/DATA1_35 ), .CK(clock), .Q(
        \U28/DATA1_35 ) );
  DFF_X2 \m2WriteBus_reg[33]  ( .D(\U3/U1/DATA1_33 ), .CK(clock), .Q(
        \U28/DATA1_33 ) );
  DFF_X2 \m2WriteAddr_reg[0]  ( .D(\eq_122/B[0] ), .CK(clock), .Q(\eq_62/B[0] ) );
  DFF_X2 \m2WriteAddr_reg[5]  ( .D(\eq_122/B[5] ), .CK(clock), .Q(\eq_62/B[5] ) );
  DFF_X2 \m2WriteAddr_reg[1]  ( .D(\eq_122/B[1] ), .CK(clock), .Q(\eq_62/B[1] ) );
  DFF_X2 \m2WriteAddr_reg[3]  ( .D(\eq_122/B[3] ), .CK(clock), .Q(\eq_62/B[3] ) );
  DFF_X2 \m2WriteAddr_reg[7]  ( .D(\eq_122/B[7] ), .CK(clock), .Q(\eq_62/B[7] ) );
  DFF_X2 \m2WriteAddr_reg[15]  ( .D(inputBaseOffset), .CK(clock), .Q(
        m2WriteAddr[15]) );
  DFF_X2 \m2WriteAddr_reg[4]  ( .D(\eq_122/B[4] ), .CK(clock), .Q(\eq_62/B[4] ) );
  DFF_X2 \m2WriteAddr_reg[2]  ( .D(\eq_122/B[2] ), .CK(clock), .Q(\eq_62/B[2] ) );
  DFF_X2 \m2WriteAddr_reg[6]  ( .D(\eq_122/B[6] ), .CK(clock), .Q(\eq_62/B[6] ) );
  DFFR_X2 \readInitial_FS_reg[5]  ( .D(\U21/Z_5 ), .CK(clock), .RN(n1531), 
        .QN(n1542) );
  DFFR_X2 m2WE_FS_reg ( .D(\U22/Z_0 ), .CK(clock), .RN(n1529), .Q(
        \U18/DATA1_0 ) );
  DFFR_X2 m2WE_FI_reg ( .D(\U25/Z_0 ), .CK(clock), .RN(n1529), .Q(
        \U22/DATA1_0 ) );
  DFFR_X2 done_FS_reg ( .D(\U23/Z_0 ), .CK(clock), .RN(n1529), .Q(
        \U19/DATA1_0 ) );
  DFFR_X2 done_FI_reg ( .D(\U26/Z_0 ), .CK(clock), .RN(n1529), .Q(
        \U23/DATA1_0 ) );
  DFFR_X2 done_Accum_reg ( .D(\U19/Z_0 ), .CK(clock), .RN(n1529), .Q(n448) );
  DFFR_X2 \readInitial_Accum_reg[4]  ( .D(\U17/Z_4 ), .CK(clock), .RN(n1531), 
        .Q(\eq_122/B[4] ) );
  DFFR_X2 \readInitial_Accum_reg[3]  ( .D(\U17/Z_3 ), .CK(clock), .RN(n1531), 
        .Q(\eq_122/B[3] ) );
  DFFR_X2 \memoryCounter_reg[2]  ( .D(n1793), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_2 ), .QN(n1726) );
  DFFR_X2 \memoryCounter_reg[12]  ( .D(n1803), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_12 ), .QN(n1771) );
  DFFR_X2 \memoryCounter_reg[8]  ( .D(n1799), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_8 ), .QN(n1752) );
  DFFR_X2 \memoryCounter_reg[10]  ( .D(n1801), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_10 ), .QN(n1761) );
  DFFR_X2 \memoryCounter_reg[6]  ( .D(n1797), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_6 ), .QN(n1744) );
  DFFR_X2 \memoryCounter_reg[4]  ( .D(n1795), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_4 ), .QN(n1735) );
  DFFR_X2 \memoryCounter_reg[13]  ( .D(n1804), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_13 ), .QN(n1775) );
  DFFR_X2 \memoryCounter_reg[1]  ( .D(n1792), .CK(clock), .RN(n1529), .Q(
        \U5/DATA1_1 ) );
  DFFR_X2 \memoryCounter_reg[11]  ( .D(n1802), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_11 ), .QN(n1717) );
  DFFR_X2 \memoryCounter_reg[9]  ( .D(n1800), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_9 ), .QN(n1715) );
  DFFR_X2 \memoryCounter_reg[7]  ( .D(n1798), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_7 ), .QN(n1716) );
  DFFR_X2 \memoryCounter_reg[5]  ( .D(n1796), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_5 ) );
  DFFR_X2 \memoryCounter_reg[3]  ( .D(n1794), .CK(clock), .RN(n1530), .Q(
        \U5/DATA1_3 ) );
  DFFR_X2 \memoryCounter_reg[14]  ( .D(n1805), .CK(clock), .RN(n1531), .Q(
        \U5/DATA1_14 ), .QN(n1784) );
  INV_X4 U3 ( .A(1'b1), .ZN(m2WriteBus[36]) );
  INV_X4 U5 ( .A(1'b1), .ZN(m2WriteBus[37]) );
  INV_X4 U7 ( .A(1'b1), .ZN(m2WriteBus[38]) );
  INV_X4 U9 ( .A(1'b1), .ZN(m2WriteBus[39]) );
  INV_X4 U12 ( .A(1'b1), .ZN(m2WriteBus[40]) );
  INV_X4 U20 ( .A(1'b1), .ZN(m2WriteBus[41]) );
  INV_X4 U22 ( .A(1'b1), .ZN(m2WriteBus[42]) );
  INV_X4 U24 ( .A(1'b1), .ZN(m2WriteBus[43]) );
  INV_X4 U28 ( .A(1'b1), .ZN(m2WriteBus[44]) );
  INV_X4 U32 ( .A(1'b1), .ZN(m2WriteBus[45]) );
  INV_X4 U36 ( .A(1'b1), .ZN(m2WriteBus[46]) );
  INV_X4 U40 ( .A(1'b1), .ZN(m2WriteBus[47]) );
  INV_X4 U44 ( .A(1'b1), .ZN(m2WriteBus[48]) );
  INV_X4 U48 ( .A(1'b1), .ZN(m2WriteBus[49]) );
  INV_X4 U52 ( .A(1'b1), .ZN(m2WriteBus[50]) );
  INV_X4 U147 ( .A(1'b1), .ZN(m2WriteBus[51]) );
  INV_X4 U149 ( .A(1'b1), .ZN(m2WriteBus[52]) );
  INV_X4 U151 ( .A(1'b1), .ZN(m2WriteBus[53]) );
  INV_X4 U153 ( .A(1'b1), .ZN(m2WriteBus[54]) );
  INV_X4 U155 ( .A(1'b1), .ZN(m2WriteBus[55]) );
  INV_X4 U157 ( .A(1'b1), .ZN(m2WriteBus[56]) );
  INV_X4 U159 ( .A(1'b1), .ZN(m2WriteBus[57]) );
  INV_X4 U161 ( .A(1'b1), .ZN(m2WriteBus[58]) );
  INV_X4 U163 ( .A(1'b1), .ZN(m2WriteBus[59]) );
  INV_X4 U165 ( .A(1'b1), .ZN(m2WriteBus[60]) );
  INV_X4 U167 ( .A(1'b1), .ZN(m2WriteBus[61]) );
  INV_X4 U169 ( .A(1'b1), .ZN(m2WriteBus[62]) );
  INV_X4 U171 ( .A(1'b1), .ZN(m2WriteBus[63]) );
  INV_X4 U173 ( .A(1'b1), .ZN(m2WriteBus[64]) );
  INV_X4 U175 ( .A(1'b1), .ZN(m2WriteBus[65]) );
  INV_X4 U177 ( .A(1'b1), .ZN(m2WriteBus[66]) );
  INV_X4 U179 ( .A(1'b1), .ZN(m2WriteBus[67]) );
  INV_X4 U181 ( .A(1'b1), .ZN(m2WriteBus[68]) );
  INV_X4 U183 ( .A(1'b1), .ZN(m2WriteBus[69]) );
  INV_X4 U185 ( .A(1'b1), .ZN(m2WriteBus[70]) );
  INV_X4 U187 ( .A(1'b1), .ZN(m2WriteBus[71]) );
  INV_X4 U189 ( .A(1'b1), .ZN(m2WriteBus[72]) );
  INV_X4 U191 ( .A(1'b1), .ZN(m2WriteBus[73]) );
  INV_X4 U193 ( .A(1'b1), .ZN(m2WriteBus[74]) );
  INV_X4 U195 ( .A(1'b1), .ZN(m2WriteBus[75]) );
  INV_X4 U197 ( .A(1'b1), .ZN(m2WriteBus[76]) );
  INV_X4 U199 ( .A(1'b1), .ZN(m2WriteBus[77]) );
  INV_X4 U201 ( .A(1'b1), .ZN(m2WriteBus[78]) );
  INV_X4 U203 ( .A(1'b1), .ZN(m2WriteBus[79]) );
  INV_X4 U205 ( .A(1'b1), .ZN(m2WriteBus[80]) );
  INV_X4 U207 ( .A(1'b1), .ZN(m2WriteBus[81]) );
  INV_X4 U209 ( .A(1'b1), .ZN(m2WriteBus[82]) );
  INV_X4 U211 ( .A(1'b1), .ZN(m2WriteBus[83]) );
  INV_X4 U213 ( .A(1'b1), .ZN(m2WriteBus[84]) );
  INV_X4 U215 ( .A(1'b1), .ZN(m2WriteBus[85]) );
  INV_X4 U217 ( .A(1'b1), .ZN(m2WriteBus[86]) );
  INV_X4 U219 ( .A(1'b1), .ZN(m2WriteBus[87]) );
  INV_X4 U221 ( .A(1'b1), .ZN(m2WriteBus[88]) );
  INV_X4 U223 ( .A(1'b1), .ZN(m2WriteBus[89]) );
  INV_X4 U225 ( .A(1'b1), .ZN(m2WriteBus[90]) );
  INV_X4 U227 ( .A(1'b1), .ZN(m2WriteBus[91]) );
  INV_X4 U229 ( .A(1'b1), .ZN(m2WriteBus[92]) );
  INV_X4 U231 ( .A(1'b1), .ZN(m2WriteBus[93]) );
  INV_X4 U233 ( .A(1'b1), .ZN(m2WriteBus[94]) );
  INV_X4 U235 ( .A(1'b1), .ZN(m2WriteBus[95]) );
  INV_X4 U237 ( .A(1'b1), .ZN(m2WriteBus[96]) );
  INV_X4 U239 ( .A(1'b1), .ZN(m2WriteBus[97]) );
  INV_X4 U241 ( .A(1'b1), .ZN(m2WriteBus[98]) );
  INV_X4 U243 ( .A(1'b1), .ZN(m2WriteBus[99]) );
  INV_X4 U245 ( .A(1'b1), .ZN(m2WriteBus[100]) );
  INV_X4 U247 ( .A(1'b1), .ZN(m2WriteBus[101]) );
  INV_X4 U249 ( .A(1'b1), .ZN(m2WriteBus[102]) );
  INV_X4 U251 ( .A(1'b1), .ZN(m2WriteBus[103]) );
  INV_X4 U253 ( .A(1'b1), .ZN(m2WriteBus[104]) );
  INV_X4 U255 ( .A(1'b1), .ZN(m2WriteBus[105]) );
  INV_X4 U257 ( .A(1'b1), .ZN(m2WriteBus[106]) );
  INV_X4 U259 ( .A(1'b1), .ZN(m2WriteBus[107]) );
  INV_X4 U261 ( .A(1'b1), .ZN(m2WriteBus[108]) );
  INV_X4 U263 ( .A(1'b1), .ZN(m2WriteBus[109]) );
  INV_X4 U265 ( .A(1'b1), .ZN(m2WriteBus[110]) );
  INV_X4 U269 ( .A(1'b1), .ZN(m2WriteBus[111]) );
  INV_X4 U273 ( .A(1'b1), .ZN(m2WriteBus[112]) );
  INV_X4 U276 ( .A(1'b1), .ZN(m2WriteBus[113]) );
  INV_X4 U281 ( .A(1'b1), .ZN(m2WriteBus[114]) );
  INV_X4 U284 ( .A(1'b1), .ZN(m2WriteBus[115]) );
  INV_X4 U287 ( .A(1'b1), .ZN(m2WriteBus[116]) );
  INV_X4 U290 ( .A(1'b1), .ZN(m2WriteBus[117]) );
  INV_X4 U292 ( .A(1'b1), .ZN(m2WriteBus[118]) );
  INV_X4 U297 ( .A(1'b1), .ZN(m2WriteBus[119]) );
  INV_X4 U301 ( .A(1'b1), .ZN(m2WriteBus[120]) );
  INV_X4 U305 ( .A(1'b1), .ZN(m2WriteBus[121]) );
  INV_X4 U308 ( .A(1'b1), .ZN(m2WriteBus[122]) );
  INV_X4 U310 ( .A(1'b1), .ZN(m2WriteBus[123]) );
  INV_X4 U314 ( .A(1'b1), .ZN(m2WriteBus[124]) );
  INV_X4 U317 ( .A(1'b1), .ZN(m2WriteBus[125]) );
  INV_X4 U320 ( .A(1'b1), .ZN(m2WriteBus[126]) );
  INV_X4 U324 ( .A(1'b1), .ZN(m2WriteBus[127]) );
  INV_X4 U327 ( .A(1'b1), .ZN(m2WriteAddr[8]) );
  INV_X4 U330 ( .A(1'b1), .ZN(m2WriteAddr[9]) );
  INV_X4 U332 ( .A(1'b1), .ZN(m2WriteAddr[10]) );
  INV_X4 U337 ( .A(1'b1), .ZN(m2WriteAddr[11]) );
  INV_X4 U342 ( .A(1'b1), .ZN(m2WriteAddr[12]) );
  INV_X4 U345 ( .A(1'b1), .ZN(m2WriteAddr[13]) );
  INV_X4 U347 ( .A(1'b1), .ZN(m2WriteAddr[14]) );
  INV_X4 U349 ( .A(1'b1), .ZN(m2ReadAddr[8]) );
  INV_X4 U351 ( .A(1'b1), .ZN(m2ReadAddr[9]) );
  INV_X4 U353 ( .A(1'b1), .ZN(m2ReadAddr[10]) );
  INV_X4 U355 ( .A(1'b1), .ZN(m2ReadAddr[11]) );
  INV_X4 U357 ( .A(1'b1), .ZN(m2ReadAddr[12]) );
  INV_X4 U359 ( .A(1'b1), .ZN(m2ReadAddr[13]) );
  INV_X4 U362 ( .A(1'b1), .ZN(m2ReadAddr[14]) );
  NAND2_X2 U364 ( .A1(n1475), .A2(n1476), .ZN(n1638) );
  NOR2_X2 U365 ( .A1(n1564), .A2(n1561), .ZN(n1486) );
  NAND2_X2 U366 ( .A1(n1705), .A2(n1704), .ZN(n1708) );
  INV_X4 U367 ( .A(n1656), .ZN(n1661) );
  OAI21_X2 U368 ( .B1(n1511), .B2(n149), .A(\U14/Z_0 ), .ZN(\U4/Z_4 ) );
  OAI21_X2 U369 ( .B1(n1512), .B2(n149), .A(\U14/Z_0 ), .ZN(\U4/Z_6 ) );
  OAI21_X2 U370 ( .B1(n1513), .B2(n149), .A(\U14/Z_0 ), .ZN(\U4/Z_5 ) );
  NOR2_X4 U371 ( .A1(\U15/DATA1_5 ), .A2(\U15/DATA1_6 ), .ZN(n1451) );
  INV_X4 U372 ( .A(n1526), .ZN(n1524) );
  NOR2_X4 U373 ( .A1(n113), .A2(n115), .ZN(n1452) );
  AND2_X4 U374 ( .A1(n1568), .A2(n1567), .ZN(n1453) );
  NOR2_X4 U375 ( .A1(n113), .A2(\U15/DATA1_5 ), .ZN(n1454) );
  AND2_X4 U376 ( .A1(n1510), .A2(n1521), .ZN(n1455) );
  OR2_X4 U377 ( .A1(n342), .A2(n343), .ZN(n1456) );
  INV_X8 U378 ( .A(n1526), .ZN(n1517) );
  INV_X4 U379 ( .A(n1516), .ZN(n1526) );
  AND2_X4 U380 ( .A1(n1722), .A2(n149), .ZN(n1459) );
  AND2_X4 U381 ( .A1(n1714), .A2(n1521), .ZN(n1460) );
  AND2_X4 U382 ( .A1(\U15/DATA1_4 ), .A2(\U15/DATA1_3 ), .ZN(n1461) );
  AND2_X4 U383 ( .A1(\U15/DATA1_5 ), .A2(n1461), .ZN(n1463) );
  OR2_X1 U384 ( .A1(n1520), .A2(\U16/DATA1_31 ), .ZN(n1464) );
  OR2_X1 U385 ( .A1(n1520), .A2(\U16/DATA1_21 ), .ZN(n1465) );
  OR2_X1 U386 ( .A1(n1520), .A2(\U16/DATA1_27 ), .ZN(n1466) );
  OR2_X1 U387 ( .A1(n1520), .A2(\U16/DATA1_25 ), .ZN(n1467) );
  OR2_X1 U388 ( .A1(n1520), .A2(\U16/DATA1_23 ), .ZN(n1468) );
  OR2_X1 U389 ( .A1(n1520), .A2(\U16/DATA1_29 ), .ZN(n1469) );
  NOR2_X1 U391 ( .A1(\U3/U1/Z_0 ), .A2(n1520), .ZN(n1471) );
  XNOR2_X1 U392 ( .A(n1690), .B(n1691), .ZN(\U16/DATA1_27 ) );
  XOR2_X1 U393 ( .A(\eq_122/B[7] ), .B(\U21/DATA1_7 ), .Z(n1548) );
  NAND2_X1 U394 ( .A1(n1493), .A2(n1702), .ZN(n1473) );
  NAND2_X2 U395 ( .A1(n1493), .A2(n1702), .ZN(n1703) );
  MUX2_X2 U396 ( .A(\U3/U1/DATA1_5 ), .B(\U3/U1/DATA2_5 ), .S(n1526), .Z(n1600) );
  INV_X2 U397 ( .A(n1486), .ZN(n1487) );
  INV_X4 U398 ( .A(n1703), .ZN(n1705) );
  XNOR2_X1 U399 ( .A(n1605), .B(n1497), .ZN(n1587) );
  NAND2_X1 U400 ( .A1(n1497), .A2(n1605), .ZN(n1593) );
  INV_X2 U401 ( .A(n1605), .ZN(n1608) );
  NAND2_X1 U402 ( .A1(\U3/U1/DATA2_16 ), .A2(n1526), .ZN(n1476) );
  INV_X4 U403 ( .A(n1569), .ZN(n1710) );
  INV_X8 U404 ( .A(n1662), .ZN(n1680) );
  NOR4_X4 U405 ( .A1(n1652), .A2(n1651), .A3(n1650), .A4(n1649), .ZN(n1654) );
  NAND3_X4 U406 ( .A1(n1681), .A2(n1680), .A3(n1679), .ZN(n1682) );
  NAND2_X2 U407 ( .A1(\U3/U1/DATA1_16 ), .A2(n1525), .ZN(n1475) );
  INV_X4 U408 ( .A(n1638), .ZN(n1644) );
  NAND2_X4 U409 ( .A1(n1661), .A2(n1660), .ZN(n1662) );
  XOR2_X1 U410 ( .A(n1644), .B(n1640), .Z(n1641) );
  XNOR2_X1 U411 ( .A(n1694), .B(n1695), .ZN(\U16/DATA1_29 ) );
  INV_X4 U412 ( .A(n1569), .ZN(n1516) );
  XOR2_X1 U413 ( .A(\eq_122/B[7] ), .B(\U17/DATA1_7 ), .Z(n1559) );
  XNOR2_X1 U414 ( .A(n1686), .B(n1687), .ZN(\U16/DATA1_25 ) );
  NAND2_X4 U415 ( .A1(n1489), .A2(n1693), .ZN(n1694) );
  XOR2_X1 U416 ( .A(\eq_122/B[3] ), .B(n1450), .Z(n1563) );
  NOR4_X4 U417 ( .A1(n1647), .A2(n1646), .A3(n1645), .A4(n1644), .ZN(n1655) );
  NOR2_X2 U418 ( .A1(n1686), .A2(n1504), .ZN(n1503) );
  NOR2_X4 U419 ( .A1(n1708), .A2(n1709), .ZN(n1712) );
  NAND3_X4 U420 ( .A1(n1653), .A2(n1654), .A3(n1655), .ZN(n1656) );
  NOR2_X4 U421 ( .A1(n1690), .A2(n1490), .ZN(n1489) );
  NOR2_X4 U427 ( .A1(n1694), .A2(n1492), .ZN(n1491) );
  NOR2_X4 U429 ( .A1(n1682), .A2(n1506), .ZN(n1505) );
  NAND2_X1 U430 ( .A1(n1707), .A2(n1483), .ZN(n1484) );
  AND2_X4 U431 ( .A1(n1700), .A2(n1699), .ZN(n1493) );
  INV_X2 U433 ( .A(n1477), .ZN(n1478) );
  NOR3_X2 U434 ( .A1(n1560), .A2(n20), .A3(n1559), .ZN(n1566) );
  NOR3_X2 U435 ( .A1(n1487), .A2(n1562), .A3(n1563), .ZN(n1565) );
  INV_X2 U436 ( .A(n1479), .ZN(n1480) );
  INV_X2 U437 ( .A(n1481), .ZN(n1482) );
  NAND3_X2 U438 ( .A1(n1453), .A2(n1566), .A3(n1565), .ZN(n1569) );
  NAND2_X1 U439 ( .A1(n1709), .A2(n1708), .ZN(n1485) );
  NAND2_X2 U440 ( .A1(n1484), .A2(n1485), .ZN(n1706) );
  INV_X1 U441 ( .A(n1708), .ZN(n1483) );
  XOR2_X2 U442 ( .A(\eq_122/B[6] ), .B(\U17/DATA1_6 ), .Z(n1562) );
  XNOR2_X1 U443 ( .A(n1698), .B(n1699), .ZN(\U16/DATA1_31 ) );
  INV_X4 U444 ( .A(n1691), .ZN(n1490) );
  INV_X4 U445 ( .A(n1695), .ZN(n1492) );
  AND2_X4 U446 ( .A1(n1653), .A2(n1648), .ZN(n1488) );
  AND2_X4 U449 ( .A1(n1680), .A2(n1666), .ZN(n1495) );
  INV_X4 U450 ( .A(n1683), .ZN(n1506) );
  INV_X4 U451 ( .A(n1687), .ZN(n1504) );
  XNOR2_X1 U452 ( .A(n1693), .B(n1489), .ZN(n1692) );
  XNOR2_X1 U453 ( .A(n1697), .B(n1491), .ZN(n1696) );
  XNOR2_X1 U454 ( .A(n1679), .B(n1673), .ZN(n1674) );
  NOR2_X1 U455 ( .A1(n1677), .A2(n1672), .ZN(n1673) );
  XNOR2_X1 U456 ( .A(n1606), .B(n1595), .ZN(n1596) );
  XNOR2_X1 U457 ( .A(n1473), .B(n1704), .ZN(\U16/DATA1_33 ) );
  XNOR2_X1 U458 ( .A(n1660), .B(n1661), .ZN(n1657) );
  XOR2_X1 U459 ( .A(n1546), .B(\eq_122/B[0] ), .Z(n1555) );
  NOR2_X1 U460 ( .A1(n1520), .A2(n1542), .ZN(\U17/Z_5 ) );
  INV_X4 U461 ( .A(n1536), .ZN(n1531) );
  INV_X4 U462 ( .A(n1536), .ZN(n1534) );
  INV_X4 U463 ( .A(n1536), .ZN(n1532) );
  INV_X4 U464 ( .A(n1536), .ZN(n1530) );
  INV_X4 U465 ( .A(n1536), .ZN(n1533) );
  INV_X4 U466 ( .A(n1536), .ZN(n1529) );
  INV_X4 U467 ( .A(n1536), .ZN(n1535) );
  INV_X4 U468 ( .A(n1455), .ZN(n1523) );
  INV_X4 U469 ( .A(rst_n), .ZN(n1536) );
  XNOR2_X2 U470 ( .A(n1682), .B(n1683), .ZN(\U16/DATA1_23 ) );
  XNOR2_X2 U471 ( .A(n1702), .B(n1493), .ZN(n1701) );
  XOR2_X2 U472 ( .A(n1689), .B(n1519), .Z(n1688) );
  XOR2_X2 U473 ( .A(n1685), .B(n1518), .Z(n1684) );
  NAND2_X2 U474 ( .A1(n1503), .A2(n1689), .ZN(n1690) );
  NAND2_X2 U475 ( .A1(n1505), .A2(n1685), .ZN(n1686) );
  NAND2_X2 U476 ( .A1(n1491), .A2(n1697), .ZN(n1698) );
  AND2_X1 U477 ( .A1(n1601), .A2(\U3/U1/Z_0 ), .ZN(n1494) );
  AND2_X1 U478 ( .A1(n1508), .A2(n1599), .ZN(n1496) );
  AND2_X1 U479 ( .A1(n1507), .A2(n1600), .ZN(n1497) );
  AND2_X1 U480 ( .A1(n1488), .A2(n1617), .ZN(n1498) );
  AND2_X1 U481 ( .A1(n1495), .A2(n1668), .ZN(n1499) );
  AND2_X1 U482 ( .A1(n1498), .A2(n1621), .ZN(n1500) );
  AND2_X1 U483 ( .A1(n1500), .A2(n1625), .ZN(n1501) );
  AND2_X1 U484 ( .A1(n1501), .A2(n1629), .ZN(n1502) );
  AND2_X1 U485 ( .A1(n1496), .A2(n1604), .ZN(n1507) );
  AND2_X1 U486 ( .A1(n1494), .A2(n1603), .ZN(n1508) );
  NAND2_X2 U487 ( .A1(n1460), .A2(n148), .ZN(n147) );
  NOR2_X2 U488 ( .A1(n342), .A2(n1807), .ZN(n319) );
  NOR2_X2 U489 ( .A1(n342), .A2(n1807), .ZN(n1522) );
  OAI21_X2 U490 ( .B1(\U15/DATA1_3 ), .B2(n149), .A(\U14/Z_0 ), .ZN(\U4/Z_3 )
         );
  INV_X4 U491 ( .A(n1528), .ZN(n1527) );
  OAI222_X2 U492 ( .A1(n285), .A2(n1812), .B1(n227), .B2(n1811), .C1(n1813), 
        .C2(n123), .ZN(n275) );
  OAI222_X2 U493 ( .A1(n276), .A2(n1812), .B1(n201), .B2(n1811), .C1(n1814), 
        .C2(n123), .ZN(n225) );
  AOI222_X1 U494 ( .A1(\U15/DATA1_3 ), .A2(n220), .B1(n237), .B2(n219), .C1(
        n238), .C2(n1835), .ZN(n236) );
  AOI222_X1 U495 ( .A1(\U15/DATA1_3 ), .A2(n213), .B1(n237), .B2(n214), .C1(
        n238), .C2(n1818), .ZN(n294) );
  AOI222_X1 U497 ( .A1(n1824), .A2(n238), .B1(n207), .B2(n237), .C1(n205), 
        .C2(\U15/DATA1_3 ), .ZN(n230) );
  AOI222_X1 U498 ( .A1(n1830), .A2(n238), .B1(n191), .B2(n237), .C1(n190), 
        .C2(\U15/DATA1_3 ), .ZN(n218) );
  AOI22_X2 U499 ( .A1(\U35/DATA1_34 ), .A2(n1452), .B1(\U35/DATA2_2 ), .B2(
        n1451), .ZN(n240) );
  AOI22_X2 U500 ( .A1(\U35/DATA1_35 ), .A2(n1452), .B1(\U35/DATA2_3 ), .B2(
        n1451), .ZN(n296) );
  AOI22_X2 U501 ( .A1(\U35/DATA1_42 ), .A2(n1452), .B1(\U35/DATA2_10 ), .B2(
        n1451), .ZN(n246) );
  AOI22_X2 U502 ( .A1(\U35/DATA1_43 ), .A2(n1452), .B1(\U35/DATA2_11 ), .B2(
        n1451), .ZN(n301) );
  AOI22_X2 U503 ( .A1(\U35/DATA1_44 ), .A2(n1452), .B1(\U35/DATA2_12 ), .B2(
        n1451), .ZN(n268) );
  AOI22_X2 U504 ( .A1(\U35/DATA1_46 ), .A2(n1452), .B1(\U35/DATA2_14 ), .B2(
        n1451), .ZN(n250) );
  AOI22_X2 U505 ( .A1(\U35/DATA1_58 ), .A2(n1452), .B1(\U35/DATA2_26 ), .B2(
        n1451), .ZN(n247) );
  AOI22_X2 U507 ( .A1(\U35/DATA1_59 ), .A2(n1452), .B1(\U35/DATA2_27 ), .B2(
        n1451), .ZN(n302) );
  AOI22_X2 U508 ( .A1(\U35/DATA1_60 ), .A2(n1452), .B1(\U35/DATA2_28 ), .B2(
        n1451), .ZN(n269) );
  AOI22_X2 U509 ( .A1(\U35/DATA1_62 ), .A2(n1452), .B1(\U35/DATA2_30 ), .B2(
        n1451), .ZN(n251) );
  XOR2_X2 U510 ( .A(n1509), .B(n1542), .Z(n1561) );
  OAI211_X2 U511 ( .C1(n344), .C2(n343), .A(n1521), .B(n345), .ZN(n342) );
  AOI21_X2 U512 ( .B1(n346), .B2(n343), .A(n1510), .ZN(n345) );
  AOI22_X2 U513 ( .A1(\U35/DATA1_41 ), .A2(n1452), .B1(\U35/DATA2_9 ), .B2(
        n1451), .ZN(n289) );
  AOI22_X2 U514 ( .A1(\U35/DATA1_45 ), .A2(n1452), .B1(\U35/DATA2_13 ), .B2(
        n1451), .ZN(n280) );
  OAI222_X2 U515 ( .A1(n123), .A2(n1815), .B1(n1811), .B2(n233), .C1(n1812), 
        .C2(n257), .ZN(n256) );
  INV_X4 U516 ( .A(n192), .ZN(n1528) );
  AOI22_X2 U517 ( .A1(n1454), .A2(\U35/DATA2_68 ), .B1(n1527), .B2(
        \U35/DATA2_36 ), .ZN(n273) );
  AOI22_X2 U518 ( .A1(\U35/DATA2_70 ), .A2(n1454), .B1(\U35/DATA2_38 ), .B2(
        n1527), .ZN(n255) );
  AOI22_X2 U519 ( .A1(\U35/DATA2_55 ), .A2(n192), .B1(\U35/DATA1_23 ), .B2(
        n1454), .ZN(n315) );
  AOI22_X2 U520 ( .A1(\U35/DATA1_55 ), .A2(n1452), .B1(\U35/DATA2_23 ), .B2(
        n1451), .ZN(n316) );
  AOI22_X2 U521 ( .A1(\U35/DATA2_50 ), .A2(n1527), .B1(\U35/DATA1_18 ), .B2(
        n1454), .ZN(n242) );
  AOI22_X2 U522 ( .A1(\U35/DATA2_51 ), .A2(n1527), .B1(\U35/DATA1_19 ), .B2(
        n1454), .ZN(n297) );
  AOI22_X2 U523 ( .A1(\U35/DATA2_52 ), .A2(n192), .B1(\U35/DATA1_20 ), .B2(
        n1454), .ZN(n270) );
  AOI22_X2 U524 ( .A1(\U35/DATA2_54 ), .A2(n192), .B1(\U35/DATA1_22 ), .B2(
        n1454), .ZN(n252) );
  AOI22_X2 U525 ( .A1(\U35/DATA1_51 ), .A2(n1452), .B1(\U35/DATA2_19 ), .B2(
        n1451), .ZN(n298) );
  AOI22_X2 U526 ( .A1(\U35/DATA1_50 ), .A2(n1452), .B1(\U35/DATA2_18 ), .B2(
        n1451), .ZN(n243) );
  AOI22_X2 U527 ( .A1(\U35/DATA1_52 ), .A2(n1452), .B1(\U35/DATA2_20 ), .B2(
        n1451), .ZN(n271) );
  AOI22_X2 U528 ( .A1(\U35/DATA1_54 ), .A2(n1452), .B1(\U35/DATA2_22 ), .B2(
        n1451), .ZN(n253) );
  AOI22_X2 U529 ( .A1(\U35/DATA1_48 ), .A2(n1452), .B1(\U35/DATA2_16 ), .B2(
        n1451), .ZN(n260) );
  AOI22_X2 U530 ( .A1(\U35/DATA1_49 ), .A2(n1452), .B1(\U35/DATA2_17 ), .B2(
        n1451), .ZN(n292) );
  AOI22_X2 U531 ( .A1(\U35/DATA1_53 ), .A2(n1452), .B1(\U35/DATA2_21 ), .B2(
        n1451), .ZN(n283) );
  AOI22_X2 U532 ( .A1(\U35/DATA2_48 ), .A2(n192), .B1(\U35/DATA1_16 ), .B2(
        n1454), .ZN(n259) );
  AOI22_X2 U533 ( .A1(\U35/DATA2_49 ), .A2(n192), .B1(\U35/DATA1_17 ), .B2(
        n1454), .ZN(n291) );
  AOI22_X2 U534 ( .A1(\U35/DATA2_53 ), .A2(n192), .B1(\U35/DATA1_21 ), .B2(
        n1454), .ZN(n282) );
  AND4_X2 U535 ( .A1(n1556), .A2(n1555), .A3(n1554), .A4(n1553), .ZN(n1510) );
  AOI21_X2 U536 ( .B1(n309), .B2(n310), .A(\U15/DATA1_3 ), .ZN(n305) );
  AOI22_X2 U537 ( .A1(\U35/DATA2_39 ), .A2(n192), .B1(\U35/DATA1_7 ), .B2(
        n1454), .ZN(n309) );
  AOI22_X2 U538 ( .A1(\U35/DATA1_39 ), .A2(n1452), .B1(\U35/DATA2_7 ), .B2(
        n1451), .ZN(n310) );
  AOI21_X2 U539 ( .B1(n307), .B2(n308), .A(n123), .ZN(n306) );
  AOI22_X2 U540 ( .A1(\U35/DATA2_47 ), .A2(n192), .B1(\U35/DATA1_15 ), .B2(
        n1454), .ZN(n307) );
  AOI22_X2 U541 ( .A1(\U35/DATA1_47 ), .A2(n1452), .B1(\U35/DATA2_15 ), .B2(
        n1451), .ZN(n308) );
  AOI21_X2 U542 ( .B1(n313), .B2(n314), .A(n123), .ZN(n312) );
  AOI22_X2 U543 ( .A1(\U35/DATA2_63 ), .A2(n192), .B1(\U35/DATA1_31 ), .B2(
        n1454), .ZN(n313) );
  AOI22_X2 U544 ( .A1(\U35/DATA1_63 ), .A2(n1452), .B1(\U35/DATA2_31 ), .B2(
        n1451), .ZN(n314) );
  OAI21_X2 U545 ( .B1(n128), .B2(n1459), .A(n1780), .ZN(n421) );
  XOR2_X2 U546 ( .A(n121), .B(\U15/DATA1_3 ), .Z(n1511) );
  XOR2_X2 U547 ( .A(n113), .B(n1463), .Z(n1512) );
  XOR2_X2 U548 ( .A(n115), .B(n1461), .Z(n1513) );
  OAI21_X2 U549 ( .B1(n311), .B2(n312), .A(\U15/DATA1_4 ), .ZN(n303) );
  OAI21_X2 U550 ( .B1(n305), .B2(n306), .A(n121), .ZN(n304) );
  AOI21_X2 U551 ( .B1(n315), .B2(n316), .A(\U15/DATA1_3 ), .ZN(n311) );
  AOI22_X2 U552 ( .A1(\U35/DATA1_40 ), .A2(n1452), .B1(\U35/DATA2_8 ), .B2(
        n1451), .ZN(n264) );
  AOI22_X2 U553 ( .A1(\U35/DATA1_56 ), .A2(n1452), .B1(\U35/DATA2_24 ), .B2(
        n1451), .ZN(n265) );
  AOI22_X2 U554 ( .A1(\U35/DATA1_57 ), .A2(n1452), .B1(\U35/DATA2_25 ), .B2(
        n1451), .ZN(n290) );
  AOI22_X2 U555 ( .A1(\U35/DATA1_61 ), .A2(n1452), .B1(\U35/DATA2_29 ), .B2(
        n1451), .ZN(n281) );
  AOI22_X2 U556 ( .A1(\U35/DATA1_32 ), .A2(n1452), .B1(\U35/DATA2_0 ), .B2(
        n1451), .ZN(n258) );
  AOI22_X2 U557 ( .A1(n1454), .A2(\U35/DATA2_65 ), .B1(n192), .B2(
        \U35/DATA2_33 ), .ZN(n293) );
  AOI22_X2 U558 ( .A1(n1454), .A2(\U35/DATA2_69 ), .B1(n1527), .B2(
        \U35/DATA2_37 ), .ZN(n284) );
  AND2_X1 U559 ( .A1(\U3/U1/DATA1_34 ), .A2(n1455), .ZN(\U20/Z_34 ) );
  INV_X4 U560 ( .A(n1520), .ZN(n1521) );
  INV_X4 U561 ( .A(start), .ZN(n1520) );
  OR2_X1 U562 ( .A1(n1520), .A2(\U16/DATA1_33 ), .ZN(n1514) );
  BUF_X4 U563 ( .A(inputBaseOffset), .Z(m2ReadAddr[15]) );
  XOR2_X1 U564 ( .A(n1676), .B(n1680), .Z(n1663) );
  NAND2_X1 U565 ( .A1(n1502), .A2(n1634), .ZN(n1639) );
  XNOR2_X1 U566 ( .A(n1600), .B(n1507), .ZN(n1584) );
  XNOR2_X1 U567 ( .A(n1601), .B(\U3/U1/Z_0 ), .ZN(n1572) );
  INV_X8 U568 ( .A(n1526), .ZN(n1525) );
  INV_X1 U569 ( .A(n1505), .ZN(n1518) );
  INV_X1 U570 ( .A(n1503), .ZN(n1519) );
  INV_X2 U571 ( .A(n1606), .ZN(n1607) );
  NOR4_X2 U580 ( .A1(n1610), .A2(n1609), .A3(n1608), .A4(n1607), .ZN(n1653) );
  XNOR2_X1 U581 ( .A(n1653), .B(n1648), .ZN(n1611) );
  XNOR2_X1 U582 ( .A(n1599), .B(n1508), .ZN(n1578) );
  NOR2_X2 U583 ( .A1(n1520), .A2(n1537), .ZN(\U21/Z_7 ) );
  NOR2_X2 U584 ( .A1(n1520), .A2(n1472), .ZN(\U17/Z_7 ) );
  XOR2_X2 U585 ( .A(n1537), .B(\eq_62/B[7] ), .Z(n1841) );
  AND2_X1 U586 ( .A1(\U18/DATA1_0 ), .A2(n1521), .ZN(\U18/Z_0 ) );
  NOR2_X2 U587 ( .A1(n1520), .A2(n1538), .ZN(\U21/Z_2 ) );
  NOR2_X2 U588 ( .A1(n1520), .A2(n1462), .ZN(\U17/Z_2 ) );
  INV_X4 U589 ( .A(n275), .ZN(n1808) );
  NOR2_X2 U592 ( .A1(n1520), .A2(n1539), .ZN(\U21/Z_1 ) );
  NOR2_X2 U593 ( .A1(n1520), .A2(n1458), .ZN(\U17/Z_1 ) );
  INV_X4 U594 ( .A(n256), .ZN(n1810) );
  NOR2_X2 U595 ( .A1(n1520), .A2(n1546), .ZN(\U21/Z_0 ) );
  NOR2_X2 U596 ( .A1(n1520), .A2(n1457), .ZN(\U17/Z_0 ) );
  NOR2_X2 U597 ( .A1(n1520), .A2(n1545), .ZN(\U21/Z_6 ) );
  NOR2_X2 U598 ( .A1(n1520), .A2(n1540), .ZN(\U17/Z_6 ) );
  INV_X4 U599 ( .A(n225), .ZN(n1809) );
  NOR2_X2 U600 ( .A1(n1520), .A2(n1541), .ZN(\U21/Z_5 ) );
  NOR2_X2 U601 ( .A1(n1520), .A2(n1543), .ZN(\U21/Z_4 ) );
  NOR2_X2 U602 ( .A1(n1520), .A2(n1481), .ZN(\U17/Z_4 ) );
  NOR2_X2 U603 ( .A1(n1520), .A2(n1544), .ZN(\U21/Z_3 ) );
  NOR2_X2 U604 ( .A1(n1520), .A2(n1474), .ZN(\U17/Z_3 ) );
  XOR2_X2 U605 ( .A(n1545), .B(\eq_122/B[6] ), .Z(n1556) );
  XOR2_X2 U606 ( .A(\eq_122/B[1] ), .B(\U21/DATA1_1 ), .Z(n1549) );
  XOR2_X2 U607 ( .A(\eq_122/B[2] ), .B(\U21/DATA1_2 ), .Z(n1547) );
  NOR3_X2 U608 ( .A1(n1549), .A2(n1548), .A3(n1547), .ZN(n1554) );
  XOR2_X2 U609 ( .A(\eq_122/B[3] ), .B(\U21/DATA1_3 ), .Z(n1552) );
  XOR2_X2 U610 ( .A(\eq_122/B[5] ), .B(\U21/DATA1_5 ), .Z(n1551) );
  XOR2_X2 U611 ( .A(\eq_122/B[4] ), .B(\U21/DATA1_4 ), .Z(n1550) );
  NOR4_X2 U612 ( .A1(n20), .A2(n1552), .A3(n1551), .A4(n1550), .ZN(n1553) );
  NAND2_X2 U613 ( .A1(\U28/DATA2_0 ), .A2(n1522), .ZN(n1557) );
  OAI221_X2 U614 ( .B1(n57), .B2(n1523), .C1(n1456), .C2(n1558), .A(n1557), 
        .ZN(\U20/Z_0 ) );
  XOR2_X2 U615 ( .A(n1457), .B(n1478), .Z(n1568) );
  XOR2_X2 U616 ( .A(n1458), .B(n1480), .Z(n1567) );
  XOR2_X2 U617 ( .A(\eq_122/B[2] ), .B(\U17/DATA1_2 ), .Z(n1560) );
  XOR2_X2 U618 ( .A(\eq_122/B[4] ), .B(n1482), .Z(n1564) );
  MUX2_X2 U619 ( .A(\U3/U1/DATA2_0 ), .B(\U3/U1/DATA1_0 ), .S(n1710), .Z(
        \U3/U1/Z_0 ) );
  NAND2_X2 U620 ( .A1(\U28/DATA2_1 ), .A2(n319), .ZN(n1570) );
  OAI221_X2 U621 ( .B1(n56), .B2(n1523), .C1(n1456), .C2(n1571), .A(n1570), 
        .ZN(\U20/Z_1 ) );
  MUX2_X2 U622 ( .A(\U3/U1/DATA2_1 ), .B(\U3/U1/DATA1_1 ), .S(n1517), .Z(n1601) );
  NOR2_X2 U623 ( .A1(n1520), .A2(n1572), .ZN(\U16/Z_1 ) );
  NAND2_X2 U624 ( .A1(\U28/DATA2_2 ), .A2(n1522), .ZN(n1573) );
  OAI221_X2 U625 ( .B1(n55), .B2(n1523), .C1(n1456), .C2(n1574), .A(n1573), 
        .ZN(\U20/Z_2 ) );
  MUX2_X2 U626 ( .A(\U3/U1/DATA2_2 ), .B(\U3/U1/DATA1_2 ), .S(n1517), .Z(n1603) );
  XNOR2_X2 U627 ( .A(n1603), .B(n1494), .ZN(n1575) );
  NOR2_X2 U628 ( .A1(n1520), .A2(n1575), .ZN(\U16/Z_2 ) );
  NAND2_X2 U629 ( .A1(\U28/DATA2_3 ), .A2(n319), .ZN(n1576) );
  OAI221_X2 U630 ( .B1(n54), .B2(n1523), .C1(n1456), .C2(n1577), .A(n1576), 
        .ZN(\U20/Z_3 ) );
  MUX2_X2 U631 ( .A(\U3/U1/DATA2_3 ), .B(\U3/U1/DATA1_3 ), .S(n1710), .Z(n1599) );
  NOR2_X2 U632 ( .A1(n1520), .A2(n1578), .ZN(\U16/Z_3 ) );
  NAND2_X2 U633 ( .A1(\U28/DATA2_4 ), .A2(n1522), .ZN(n1579) );
  OAI221_X2 U634 ( .B1(n53), .B2(n1523), .C1(n1456), .C2(n1580), .A(n1579), 
        .ZN(\U20/Z_4 ) );
  MUX2_X2 U635 ( .A(\U3/U1/DATA2_4 ), .B(\U3/U1/DATA1_4 ), .S(n1517), .Z(n1604) );
  XNOR2_X2 U636 ( .A(n1604), .B(n1496), .ZN(n1581) );
  NOR2_X2 U637 ( .A1(n1520), .A2(n1581), .ZN(\U16/Z_4 ) );
  NAND2_X2 U638 ( .A1(\U28/DATA2_5 ), .A2(n319), .ZN(n1582) );
  OAI221_X2 U639 ( .B1(n52), .B2(n1523), .C1(n1456), .C2(n1583), .A(n1582), 
        .ZN(\U20/Z_5 ) );
  NOR2_X2 U640 ( .A1(n1520), .A2(n1584), .ZN(\U16/Z_5 ) );
  NAND2_X2 U641 ( .A1(\U28/DATA2_6 ), .A2(n1522), .ZN(n1585) );
  OAI221_X2 U642 ( .B1(n51), .B2(n1523), .C1(n1456), .C2(n1586), .A(n1585), 
        .ZN(\U20/Z_6 ) );
  MUX2_X2 U643 ( .A(\U3/U1/DATA2_6 ), .B(\U3/U1/DATA1_6 ), .S(n1525), .Z(n1605) );
  NOR2_X2 U644 ( .A1(n1520), .A2(n1587), .ZN(\U16/Z_6 ) );
  NAND2_X2 U645 ( .A1(\U28/DATA2_7 ), .A2(n319), .ZN(n1588) );
  OAI221_X2 U646 ( .B1(n50), .B2(n1523), .C1(n1456), .C2(n1589), .A(n1588), 
        .ZN(\U20/Z_7 ) );
  MUX2_X2 U647 ( .A(\U3/U1/DATA2_7 ), .B(\U3/U1/DATA1_7 ), .S(n1517), .Z(n1602) );
  INV_X4 U648 ( .A(n1602), .ZN(n1594) );
  XNOR2_X2 U649 ( .A(n1594), .B(n1593), .ZN(n1590) );
  NOR2_X2 U650 ( .A1(n1520), .A2(n1590), .ZN(\U16/Z_7 ) );
  NAND2_X2 U651 ( .A1(\U28/DATA2_8 ), .A2(n1522), .ZN(n1591) );
  OAI221_X2 U652 ( .B1(n49), .B2(n1523), .C1(n1456), .C2(n1592), .A(n1591), 
        .ZN(\U20/Z_8 ) );
  MUX2_X2 U653 ( .A(\U3/U1/DATA2_8 ), .B(\U3/U1/DATA1_8 ), .S(n1525), .Z(n1606) );
  NOR2_X2 U654 ( .A1(n1594), .A2(n1593), .ZN(n1595) );
  NOR2_X2 U655 ( .A1(n1520), .A2(n1596), .ZN(\U16/Z_8 ) );
  NAND2_X2 U656 ( .A1(\U28/DATA2_9 ), .A2(n319), .ZN(n1597) );
  OAI221_X2 U657 ( .B1(n48), .B2(n1523), .C1(n1456), .C2(n1598), .A(n1597), 
        .ZN(\U20/Z_9 ) );
  NAND4_X2 U658 ( .A1(n1601), .A2(n1600), .A3(\U3/U1/Z_0 ), .A4(n1599), .ZN(
        n1610) );
  NAND3_X2 U659 ( .A1(n1604), .A2(n1603), .A3(n1602), .ZN(n1609) );
  MUX2_X2 U660 ( .A(\U3/U1/DATA2_9 ), .B(\U3/U1/DATA1_9 ), .S(n1525), .Z(n1648) );
  NOR2_X2 U661 ( .A1(n1520), .A2(n1611), .ZN(\U16/Z_9 ) );
  NAND2_X2 U662 ( .A1(\U28/DATA2_10 ), .A2(n1522), .ZN(n1612) );
  OAI221_X2 U663 ( .B1(n47), .B2(n1523), .C1(n1456), .C2(n1613), .A(n1612), 
        .ZN(\U20/Z_10 ) );
  MUX2_X2 U664 ( .A(\U3/U1/DATA2_10 ), .B(\U3/U1/DATA1_10 ), .S(n1525), .Z(
        n1617) );
  INV_X4 U665 ( .A(n1617), .ZN(n1647) );
  XOR2_X2 U666 ( .A(n1647), .B(n1488), .Z(n1614) );
  NOR2_X2 U667 ( .A1(n1520), .A2(n1614), .ZN(\U16/Z_10 ) );
  NAND2_X2 U668 ( .A1(\U28/DATA2_11 ), .A2(n319), .ZN(n1615) );
  OAI221_X2 U669 ( .B1(n46), .B2(n1523), .C1(n1456), .C2(n1616), .A(n1615), 
        .ZN(\U20/Z_11 ) );
  MUX2_X2 U670 ( .A(\U3/U1/DATA2_11 ), .B(\U3/U1/DATA1_11 ), .S(n1525), .Z(
        n1621) );
  INV_X4 U671 ( .A(n1621), .ZN(n1651) );
  XOR2_X2 U672 ( .A(n1651), .B(n1498), .Z(n1618) );
  NOR2_X2 U673 ( .A1(n1520), .A2(n1618), .ZN(\U16/Z_11 ) );
  NAND2_X2 U674 ( .A1(\U28/DATA2_12 ), .A2(n1522), .ZN(n1619) );
  OAI221_X2 U675 ( .B1(n45), .B2(n1523), .C1(n1456), .C2(n1620), .A(n1619), 
        .ZN(\U20/Z_12 ) );
  MUX2_X2 U676 ( .A(\U3/U1/DATA2_12 ), .B(\U3/U1/DATA1_12 ), .S(n1525), .Z(
        n1625) );
  INV_X4 U677 ( .A(n1625), .ZN(n1646) );
  XOR2_X2 U678 ( .A(n1646), .B(n1500), .Z(n1622) );
  NOR2_X2 U679 ( .A1(n1520), .A2(n1622), .ZN(\U16/Z_12 ) );
  NAND2_X2 U680 ( .A1(\U28/DATA2_13 ), .A2(n319), .ZN(n1623) );
  OAI221_X2 U681 ( .B1(n44), .B2(n1523), .C1(n1456), .C2(n1624), .A(n1623), 
        .ZN(\U20/Z_13 ) );
  MUX2_X2 U682 ( .A(\U3/U1/DATA2_13 ), .B(\U3/U1/DATA1_13 ), .S(n1525), .Z(
        n1629) );
  INV_X4 U683 ( .A(n1629), .ZN(n1650) );
  XOR2_X2 U684 ( .A(n1650), .B(n1501), .Z(n1626) );
  NOR2_X2 U685 ( .A1(n1520), .A2(n1626), .ZN(\U16/Z_13 ) );
  NAND2_X2 U686 ( .A1(\U28/DATA2_14 ), .A2(n1522), .ZN(n1627) );
  OAI221_X2 U687 ( .B1(n42), .B2(n1523), .C1(n1456), .C2(n1628), .A(n1627), 
        .ZN(\U20/Z_14 ) );
  MUX2_X2 U688 ( .A(\U3/U1/DATA2_14 ), .B(\U3/U1/DATA1_14 ), .S(n1525), .Z(
        n1634) );
  INV_X4 U689 ( .A(n1634), .ZN(n1645) );
  XOR2_X2 U690 ( .A(n1645), .B(n1502), .Z(n1630) );
  NOR2_X2 U691 ( .A1(n1520), .A2(n1630), .ZN(\U16/Z_14 ) );
  NAND2_X2 U692 ( .A1(\U28/DATA2_15 ), .A2(n319), .ZN(n1631) );
  OAI221_X2 U693 ( .B1(n41), .B2(n1523), .C1(n1456), .C2(n1632), .A(n1631), 
        .ZN(\U20/Z_15 ) );
  MUX2_X2 U694 ( .A(\U3/U1/DATA2_15 ), .B(\U3/U1/DATA1_15 ), .S(n1525), .Z(
        n1633) );
  INV_X4 U695 ( .A(n1633), .ZN(n1649) );
  XNOR2_X2 U696 ( .A(n1649), .B(n1639), .ZN(n1635) );
  NOR2_X2 U697 ( .A1(n1520), .A2(n1635), .ZN(\U16/Z_15 ) );
  NAND2_X2 U698 ( .A1(\U28/DATA2_16 ), .A2(n1522), .ZN(n1636) );
  OAI221_X2 U699 ( .B1(n40), .B2(n1523), .C1(n1456), .C2(n1637), .A(n1636), 
        .ZN(\U20/Z_16 ) );
  NOR2_X2 U700 ( .A1(n1649), .A2(n1639), .ZN(n1640) );
  NOR2_X2 U701 ( .A1(n1520), .A2(n1641), .ZN(\U16/Z_16 ) );
  NAND2_X2 U702 ( .A1(\U28/DATA2_17 ), .A2(n319), .ZN(n1642) );
  OAI221_X2 U703 ( .B1(n39), .B2(n1523), .C1(n1456), .C2(n1643), .A(n1642), 
        .ZN(\U20/Z_17 ) );
  MUX2_X2 U704 ( .A(\U3/U1/DATA2_17 ), .B(\U3/U1/DATA1_17 ), .S(n1524), .Z(
        n1660) );
  INV_X4 U705 ( .A(n1648), .ZN(n1652) );
  NOR2_X2 U706 ( .A1(n1520), .A2(n1657), .ZN(\U16/Z_17 ) );
  NAND2_X2 U707 ( .A1(\U28/DATA2_18 ), .A2(n1522), .ZN(n1658) );
  OAI221_X2 U708 ( .B1(n38), .B2(n1523), .C1(n1456), .C2(n1659), .A(n1658), 
        .ZN(\U20/Z_18 ) );
  MUX2_X2 U709 ( .A(\U3/U1/DATA2_18 ), .B(\U3/U1/DATA1_18 ), .S(n1525), .Z(
        n1666) );
  INV_X4 U710 ( .A(n1666), .ZN(n1676) );
  NOR2_X2 U711 ( .A1(n1520), .A2(n1663), .ZN(\U16/Z_18 ) );
  NAND2_X2 U712 ( .A1(\U28/DATA2_19 ), .A2(n319), .ZN(n1664) );
  OAI221_X2 U713 ( .B1(n37), .B2(n1523), .C1(n1456), .C2(n1665), .A(n1664), 
        .ZN(\U20/Z_19 ) );
  MUX2_X2 U714 ( .A(\U3/U1/DATA2_19 ), .B(\U3/U1/DATA1_19 ), .S(n1524), .Z(
        n1668) );
  INV_X4 U715 ( .A(n1668), .ZN(n1678) );
  XOR2_X2 U716 ( .A(n1678), .B(n1495), .Z(n1667) );
  NOR2_X2 U717 ( .A1(n1520), .A2(n1667), .ZN(\U16/Z_19 ) );
  NOR2_X2 U718 ( .A1(n36), .A2(n1523), .ZN(\U20/Z_20 ) );
  MUX2_X2 U719 ( .A(\U3/U1/DATA2_20 ), .B(\U3/U1/DATA1_20 ), .S(n1525), .Z(
        n1670) );
  INV_X4 U720 ( .A(n1670), .ZN(n1675) );
  XOR2_X2 U721 ( .A(n1675), .B(n1499), .Z(n1669) );
  NOR2_X2 U722 ( .A1(n1520), .A2(n1669), .ZN(\U16/Z_20 ) );
  NAND2_X2 U723 ( .A1(n35), .A2(n1455), .ZN(\U20/Z_21 ) );
  NAND2_X2 U724 ( .A1(n1499), .A2(n1670), .ZN(n1672) );
  MUX2_X2 U725 ( .A(\U3/U1/DATA2_21 ), .B(\U3/U1/DATA1_21 ), .S(n1524), .Z(
        n1671) );
  INV_X4 U726 ( .A(n1671), .ZN(n1677) );
  XOR2_X2 U727 ( .A(n1672), .B(n1677), .Z(\U16/DATA1_21 ) );
  NOR2_X2 U728 ( .A1(n34), .A2(n1523), .ZN(\U20/Z_22 ) );
  MUX2_X2 U729 ( .A(\U3/U1/DATA2_22 ), .B(\U3/U1/DATA1_22 ), .S(n1524), .Z(
        n1679) );
  NOR2_X2 U730 ( .A1(n1520), .A2(n1674), .ZN(\U16/Z_22 ) );
  NAND2_X2 U731 ( .A1(n33), .A2(n1455), .ZN(\U20/Z_23 ) );
  NOR4_X2 U732 ( .A1(n1678), .A2(n1677), .A3(n1676), .A4(n1675), .ZN(n1681) );
  MUX2_X2 U733 ( .A(\U3/U1/DATA2_23 ), .B(\U3/U1/DATA1_23 ), .S(n1524), .Z(
        n1683) );
  NOR2_X2 U734 ( .A1(n32), .A2(n1523), .ZN(\U20/Z_24 ) );
  MUX2_X2 U735 ( .A(\U3/U1/DATA2_24 ), .B(\U3/U1/DATA1_24 ), .S(n1524), .Z(
        n1685) );
  NOR2_X2 U736 ( .A1(n1520), .A2(n1684), .ZN(\U16/Z_24 ) );
  NAND2_X2 U737 ( .A1(n31), .A2(n1455), .ZN(\U20/Z_25 ) );
  MUX2_X2 U738 ( .A(\U3/U1/DATA2_25 ), .B(\U3/U1/DATA1_25 ), .S(n1524), .Z(
        n1687) );
  NOR2_X2 U739 ( .A1(n30), .A2(n1523), .ZN(\U20/Z_26 ) );
  MUX2_X2 U740 ( .A(\U3/U1/DATA2_26 ), .B(\U3/U1/DATA1_26 ), .S(n1524), .Z(
        n1689) );
  NOR2_X2 U741 ( .A1(n1520), .A2(n1688), .ZN(\U16/Z_26 ) );
  NAND2_X2 U742 ( .A1(n29), .A2(n1455), .ZN(\U20/Z_27 ) );
  MUX2_X2 U743 ( .A(\U3/U1/DATA2_27 ), .B(\U3/U1/DATA1_27 ), .S(n1524), .Z(
        n1691) );
  NOR2_X2 U744 ( .A1(n28), .A2(n1523), .ZN(\U20/Z_28 ) );
  MUX2_X2 U745 ( .A(\U3/U1/DATA2_28 ), .B(\U3/U1/DATA1_28 ), .S(n1524), .Z(
        n1693) );
  NOR2_X2 U746 ( .A1(n1520), .A2(n1692), .ZN(\U16/Z_28 ) );
  NAND2_X2 U747 ( .A1(n27), .A2(n1455), .ZN(\U20/Z_29 ) );
  MUX2_X2 U748 ( .A(\U3/U1/DATA2_29 ), .B(\U3/U1/DATA1_29 ), .S(n1524), .Z(
        n1695) );
  NOR2_X2 U749 ( .A1(n26), .A2(n1523), .ZN(\U20/Z_30 ) );
  MUX2_X2 U750 ( .A(\U3/U1/DATA2_30 ), .B(\U3/U1/DATA1_30 ), .S(n1524), .Z(
        n1697) );
  NOR2_X2 U751 ( .A1(n1520), .A2(n1696), .ZN(\U16/Z_30 ) );
  NAND2_X2 U752 ( .A1(n25), .A2(n1455), .ZN(\U20/Z_31 ) );
  MUX2_X2 U753 ( .A(\U3/U1/DATA2_31 ), .B(\U3/U1/DATA1_31 ), .S(n1524), .Z(
        n1699) );
  NOR2_X2 U754 ( .A1(n24), .A2(n1523), .ZN(\U20/Z_32 ) );
  MUX2_X2 U755 ( .A(\U3/U1/DATA2_32 ), .B(\U3/U1/DATA1_32 ), .S(n1524), .Z(
        n1702) );
  INV_X4 U756 ( .A(n1698), .ZN(n1700) );
  NOR2_X2 U757 ( .A1(n1520), .A2(n1701), .ZN(\U16/Z_32 ) );
  NAND2_X2 U758 ( .A1(n23), .A2(n1455), .ZN(\U20/Z_33 ) );
  MUX2_X2 U759 ( .A(\U3/U1/DATA2_33 ), .B(\U3/U1/DATA1_33 ), .S(n1524), .Z(
        n1704) );
  MUX2_X2 U760 ( .A(\U3/U1/DATA2_34 ), .B(\U3/U1/DATA1_34 ), .S(n1524), .Z(
        n1707) );
  NOR2_X2 U761 ( .A1(n1520), .A2(n1706), .ZN(\U16/Z_34 ) );
  NAND2_X2 U762 ( .A1(n21), .A2(n1455), .ZN(\U20/Z_35 ) );
  INV_X4 U763 ( .A(n1707), .ZN(n1709) );
  MUX2_X2 U764 ( .A(\U3/U1/DATA2_35 ), .B(\U3/U1/DATA1_35 ), .S(n1524), .Z(
        n1711) );
  XNOR2_X2 U765 ( .A(n1712), .B(n1711), .ZN(n1713) );
  NAND2_X2 U766 ( .A1(n1521), .A2(n1713), .ZN(\U16/Z_35 ) );
  NAND2_X2 U767 ( .A1(n208), .A2(n1452), .ZN(n1721) );
  INV_X4 U768 ( .A(n1721), .ZN(n1714) );
  NAND3_X2 U769 ( .A1(\U5/DATA1_1 ), .A2(\U5/DATA1_0 ), .A3(\U5/DATA1_2 ), 
        .ZN(n1729) );
  INV_X4 U770 ( .A(n1729), .ZN(n1732) );
  NAND3_X2 U771 ( .A1(\U5/DATA1_4 ), .A2(\U5/DATA1_3 ), .A3(n1732), .ZN(n1738)
         );
  INV_X4 U772 ( .A(n1738), .ZN(n1741) );
  NAND3_X2 U773 ( .A1(\U5/DATA1_6 ), .A2(\U5/DATA1_5 ), .A3(n1741), .ZN(n1747)
         );
  INV_X4 U774 ( .A(n1747), .ZN(n1755) );
  NOR3_X2 U775 ( .A1(n1717), .A2(n1716), .A3(n1715), .ZN(n1719) );
  NOR4_X2 U776 ( .A1(\U5/DATA1_10 ), .A2(\U5/DATA1_8 ), .A3(\U5/DATA1_13 ), 
        .A4(\U5/DATA1_12 ), .ZN(n1718) );
  NAND4_X2 U777 ( .A1(\U5/DATA1_14 ), .A2(n1755), .A3(n1719), .A4(n1718), .ZN(
        n148) );
  NOR2_X2 U778 ( .A1(n147), .A2(n128), .ZN(n1723) );
  INV_X4 U779 ( .A(n148), .ZN(n1720) );
  NAND2_X2 U780 ( .A1(n1460), .A2(n1720), .ZN(n1722) );
  NAND2_X2 U781 ( .A1(n1721), .A2(n1521), .ZN(n149) );
  INV_X4 U782 ( .A(n147), .ZN(n1765) );
  NAND2_X2 U783 ( .A1(n1765), .A2(n128), .ZN(n1780) );
  NAND2_X2 U784 ( .A1(n1459), .A2(n1780), .ZN(n1725) );
  MUX2_X2 U785 ( .A(n1723), .B(n1725), .S(\U5/DATA1_1 ), .Z(n1792) );
  NAND2_X2 U786 ( .A1(\U5/DATA1_0 ), .A2(n1726), .ZN(n1724) );
  MUX2_X2 U787 ( .A(n1726), .B(n1724), .S(\U5/DATA1_1 ), .Z(n1728) );
  INV_X4 U788 ( .A(n1725), .ZN(n1727) );
  OAI22_X2 U789 ( .A1(n147), .A2(n1728), .B1(n1727), .B2(n1726), .ZN(n1793) );
  NOR2_X2 U790 ( .A1(n147), .A2(n1729), .ZN(n1731) );
  NAND2_X2 U791 ( .A1(n1729), .A2(n1765), .ZN(n1730) );
  NAND2_X2 U792 ( .A1(n1459), .A2(n1730), .ZN(n1734) );
  MUX2_X2 U793 ( .A(n1731), .B(n1734), .S(\U5/DATA1_3 ), .Z(n1794) );
  NAND2_X2 U794 ( .A1(n1732), .A2(n1735), .ZN(n1733) );
  MUX2_X2 U795 ( .A(n1735), .B(n1733), .S(\U5/DATA1_3 ), .Z(n1737) );
  INV_X4 U796 ( .A(n1734), .ZN(n1736) );
  OAI22_X2 U797 ( .A1(n147), .A2(n1737), .B1(n1736), .B2(n1735), .ZN(n1795) );
  NOR2_X2 U798 ( .A1(n147), .A2(n1738), .ZN(n1740) );
  NAND2_X2 U799 ( .A1(n1738), .A2(n1765), .ZN(n1739) );
  NAND2_X2 U800 ( .A1(n1459), .A2(n1739), .ZN(n1743) );
  MUX2_X2 U801 ( .A(n1740), .B(n1743), .S(\U5/DATA1_5 ), .Z(n1796) );
  NAND2_X2 U802 ( .A1(n1741), .A2(n1744), .ZN(n1742) );
  MUX2_X2 U803 ( .A(n1744), .B(n1742), .S(\U5/DATA1_5 ), .Z(n1746) );
  INV_X4 U804 ( .A(n1743), .ZN(n1745) );
  OAI22_X2 U805 ( .A1(n147), .A2(n1746), .B1(n1745), .B2(n1744), .ZN(n1797) );
  NOR2_X2 U806 ( .A1(n147), .A2(n1747), .ZN(n1749) );
  NAND2_X2 U807 ( .A1(n1747), .A2(n1765), .ZN(n1748) );
  NAND2_X2 U808 ( .A1(n1459), .A2(n1748), .ZN(n1751) );
  MUX2_X2 U809 ( .A(n1749), .B(n1751), .S(\U5/DATA1_7 ), .Z(n1798) );
  NAND2_X2 U810 ( .A1(n1755), .A2(n1752), .ZN(n1750) );
  MUX2_X2 U811 ( .A(n1752), .B(n1750), .S(\U5/DATA1_7 ), .Z(n1754) );
  INV_X4 U812 ( .A(n1751), .ZN(n1753) );
  OAI22_X2 U813 ( .A1(n147), .A2(n1754), .B1(n1753), .B2(n1752), .ZN(n1799) );
  NAND3_X2 U814 ( .A1(\U5/DATA1_8 ), .A2(\U5/DATA1_7 ), .A3(n1755), .ZN(n1758)
         );
  NOR2_X2 U815 ( .A1(n147), .A2(n1758), .ZN(n1757) );
  NAND2_X2 U816 ( .A1(n1758), .A2(n1765), .ZN(n1756) );
  NAND2_X2 U817 ( .A1(n1459), .A2(n1756), .ZN(n1760) );
  MUX2_X2 U818 ( .A(n1757), .B(n1760), .S(\U5/DATA1_9 ), .Z(n1800) );
  INV_X4 U819 ( .A(n1758), .ZN(n1764) );
  NAND2_X2 U820 ( .A1(n1764), .A2(n1761), .ZN(n1759) );
  MUX2_X2 U821 ( .A(n1761), .B(n1759), .S(\U5/DATA1_9 ), .Z(n1763) );
  INV_X4 U822 ( .A(n1760), .ZN(n1762) );
  OAI22_X2 U823 ( .A1(n147), .A2(n1763), .B1(n1762), .B2(n1761), .ZN(n1801) );
  NAND3_X2 U824 ( .A1(\U5/DATA1_10 ), .A2(\U5/DATA1_9 ), .A3(n1764), .ZN(n1768) );
  NOR2_X2 U825 ( .A1(n147), .A2(n1768), .ZN(n1767) );
  NAND2_X2 U826 ( .A1(n1768), .A2(n1765), .ZN(n1766) );
  NAND2_X2 U827 ( .A1(n1459), .A2(n1766), .ZN(n1770) );
  MUX2_X2 U828 ( .A(n1767), .B(n1770), .S(\U5/DATA1_11 ), .Z(n1802) );
  INV_X4 U829 ( .A(n1768), .ZN(n1774) );
  NAND2_X2 U830 ( .A1(n1774), .A2(n1771), .ZN(n1769) );
  MUX2_X2 U831 ( .A(n1771), .B(n1769), .S(\U5/DATA1_11 ), .Z(n1773) );
  INV_X4 U832 ( .A(n1770), .ZN(n1772) );
  OAI22_X2 U833 ( .A1(n147), .A2(n1773), .B1(n1772), .B2(n1771), .ZN(n1803) );
  NAND3_X2 U834 ( .A1(\U5/DATA1_12 ), .A2(\U5/DATA1_11 ), .A3(n1774), .ZN(
        n1777) );
  XOR2_X2 U835 ( .A(n1777), .B(\U5/DATA1_13 ), .Z(n1776) );
  OAI22_X2 U836 ( .A1(n147), .A2(n1776), .B1(n1459), .B2(n1775), .ZN(n1804) );
  INV_X4 U837 ( .A(n1777), .ZN(n1778) );
  NAND2_X2 U838 ( .A1(\U5/DATA1_13 ), .A2(n1778), .ZN(n1785) );
  XOR2_X2 U839 ( .A(n1785), .B(\U5/DATA1_14 ), .Z(n1779) );
  OAI22_X2 U840 ( .A1(n147), .A2(n1779), .B1(n1459), .B2(n1784), .ZN(n1805) );
  INV_X4 U841 ( .A(n1785), .ZN(n1781) );
  NAND2_X2 U842 ( .A1(n1781), .A2(\U5/DATA1_14 ), .ZN(n1782) );
  NAND2_X2 U843 ( .A1(n1460), .A2(n1782), .ZN(n1783) );
  NAND2_X2 U844 ( .A1(n1459), .A2(n1783), .ZN(n1787) );
  NOR3_X2 U845 ( .A1(n1785), .A2(n147), .A3(n1784), .ZN(n1786) );
  MUX2_X2 U846 ( .A(n1787), .B(n1786), .S(n127), .Z(n420) );
  NAND4_X2 U847 ( .A1(n1791), .A2(n1790), .A3(n1789), .A4(n1788), .ZN(n371) );
  NAND4_X2 U848 ( .A1(\U28/DATA1_23 ), .A2(\U28/DATA1_21 ), .A3(\U28/DATA1_27 ), .A4(\U28/DATA1_25 ), .ZN(n372) );
  XOR2_X2 U849 ( .A(\eq_62/B[3] ), .B(\U21/DATA1_3 ), .Z(n358) );
  XOR2_X2 U850 ( .A(\eq_62/B[4] ), .B(\U21/DATA1_4 ), .Z(n359) );
  XOR2_X2 U851 ( .A(\eq_62/B[5] ), .B(\U21/DATA1_5 ), .Z(n360) );
  XOR2_X2 U852 ( .A(\eq_62/B[6] ), .B(\U21/DATA1_6 ), .Z(n361) );
  XOR2_X2 U853 ( .A(\eq_62/B[0] ), .B(\U21/DATA1_0 ), .Z(n355) );
  XOR2_X2 U854 ( .A(\eq_62/B[1] ), .B(\U21/DATA1_1 ), .Z(n356) );
  XOR2_X2 U855 ( .A(\eq_62/B[2] ), .B(\U21/DATA1_2 ), .Z(n357) );
  INV_X4 U856 ( .A(n343), .ZN(n1807) );
  INV_X4 U857 ( .A(\U14/Z_0 ), .ZN(n1806) );
  INV_X4 U858 ( .A(n237), .ZN(n1811) );
  INV_X4 U859 ( .A(n238), .ZN(n1812) );
  INV_X4 U860 ( .A(n286), .ZN(n1813) );
  INV_X4 U861 ( .A(n277), .ZN(n1814) );
  INV_X4 U862 ( .A(n261), .ZN(n1815) );
  INV_X4 U863 ( .A(n302), .ZN(n1816) );
  INV_X4 U864 ( .A(n301), .ZN(n1817) );
  INV_X4 U865 ( .A(n295), .ZN(n1818) );
  INV_X4 U866 ( .A(n296), .ZN(n1819) );
  INV_X4 U867 ( .A(n290), .ZN(n1820) );
  INV_X4 U868 ( .A(n289), .ZN(n1821) );
  INV_X4 U869 ( .A(n281), .ZN(n1822) );
  INV_X4 U870 ( .A(n280), .ZN(n1823) );
  INV_X4 U871 ( .A(n272), .ZN(n1824) );
  INV_X4 U872 ( .A(n269), .ZN(n1825) );
  INV_X4 U873 ( .A(n268), .ZN(n1826) );
  INV_X4 U874 ( .A(n265), .ZN(n1827) );
  INV_X4 U875 ( .A(n264), .ZN(n1828) );
  INV_X4 U876 ( .A(n258), .ZN(n1829) );
  INV_X4 U877 ( .A(n254), .ZN(n1830) );
  INV_X4 U878 ( .A(n251), .ZN(n1831) );
  INV_X4 U879 ( .A(n250), .ZN(n1832) );
  INV_X4 U880 ( .A(n247), .ZN(n1833) );
  INV_X4 U881 ( .A(n246), .ZN(n1834) );
  INV_X4 U882 ( .A(n239), .ZN(n1835) );
  INV_X4 U883 ( .A(n240), .ZN(n1836) );
  INV_X4 U884 ( .A(n293), .ZN(n1837) );
  INV_X4 U885 ( .A(n284), .ZN(n1838) );
  INV_X4 U886 ( .A(n273), .ZN(n1839) );
  INV_X4 U887 ( .A(n255), .ZN(n1840) );
  NAND3_X2 U888 ( .A1(n353), .A2(n354), .A3(n1841), .ZN(n343) );
endmodule


module Cdf_Fetch ( clock, reset_n, start, ReadBus, ReadAddr, AccumlateOut, 
        StartOut, StoreAddress, input_base_offset, done );
  input [35:0] ReadBus;
  output [15:0] ReadAddr;
  output [19:0] AccumlateOut;
  output [15:0] StoreAddress;
  input clock, reset_n, start, input_base_offset;
  output StartOut, done;
  wire   \U3/U1/DATA1_1 , \U3/U1/DATA1_2 , \U3/U1/DATA1_3 , \U3/U1/DATA1_4 ,
         \U3/U1/DATA1_5 , \U3/U1/DATA1_6 , \U3/U1/DATA1_7 , \U11/DATA1_0 ,
         \U11/DATA1_1 , \U11/DATA1_2 , \U11/DATA1_3 , \U11/DATA1_4 ,
         \U11/DATA1_5 , \U11/DATA1_6 , \U11/DATA1_7 , \U11/DATA1_8 ,
         \U11/DATA1_9 , \U11/DATA1_10 , \U11/DATA1_11 , \U11/DATA1_12 ,
         \U11/DATA1_13 , \U11/DATA1_14 , \U11/DATA1_15 , \U11/DATA1_16 ,
         \U11/DATA1_17 , \U11/DATA1_18 , \U11/DATA1_19 , \U10/Z_0 , \U10/Z_1 ,
         \U10/Z_2 , \U10/Z_3 , \U10/Z_4 , \U10/Z_5 , \U10/Z_6 , \U10/Z_7 ,
         \U10/Z_8 , \U10/Z_9 , \U10/Z_10 , \U10/Z_11 , \U10/Z_12 , \U10/Z_13 ,
         \U10/Z_14 , \U10/Z_15 , \U10/DATA1_0 , \U10/DATA1_1 , \U10/DATA1_2 ,
         \U10/DATA1_3 , \U10/DATA1_4 , \U10/DATA1_5 , \U10/DATA1_6 ,
         \U10/DATA1_7 , \U10/DATA1_8 , \U10/DATA1_9 , \U10/DATA1_10 ,
         \U10/DATA1_11 , \U10/DATA1_12 , \U10/DATA1_13 , \U10/DATA1_14 ,
         \U10/DATA1_15 , \U9/Z_0 , \U9/DATA1_0 , \U8/Z_0 , \U8/DATA1_0 ,
         \U7/Z_0 , \U7/Z_1 , \U7/Z_2 , \U7/Z_3 , \U7/Z_4 , \U7/Z_5 , \U7/Z_6 ,
         \U7/Z_7 , \U7/Z_8 , \U7/Z_9 , \U7/Z_10 , \U7/Z_11 , \U7/Z_12 ,
         \U7/Z_13 , \U7/Z_14 , \U7/Z_15 , \U7/Z_16 , \U7/Z_17 , \U7/Z_18 ,
         \U7/Z_19 , \U5/Z_0 , \U5/Z_1 , \U5/Z_2 , \U5/Z_3 , \U5/Z_4 , \U5/Z_5 ,
         \U5/Z_6 , \U5/Z_7 , \U5/Z_8 , \U5/Z_9 , \U5/Z_10 , \U5/Z_11 ,
         \U5/Z_12 , \U5/Z_13 , \U5/Z_14 , \U5/DATA1_1 , \U5/DATA1_2 ,
         \U5/DATA1_3 , \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 , \U5/DATA1_7 ,
         \U5/DATA1_8 , \U5/DATA1_9 , \U5/DATA1_10 , \U5/DATA1_11 ,
         \U5/DATA1_12 , \U5/DATA1_13 , \U5/DATA1_14 , \U4/Z_0 , \U4/CONTROL2 ,
         \U4/DATA3_0 , \add_69/carry[8] , \add_69/carry[7] , \add_69/carry[6] ,
         \add_69/carry[5] , \add_69/carry[4] , \add_69/carry[3] ,
         \add_69/carry[2] , \add_69/A[0] , \add_69/A[1] , \add_69/A[2] ,
         \add_69/A[3] , \add_69/A[4] , \add_69/A[5] , \add_69/A[6] ,
         \add_69/A[7] , \add_69/A[8] , \add_66/carry[15] , \add_66/carry[14] ,
         \add_66/carry[12] , \add_66/carry[11] , \add_66/carry[10] ,
         \add_66/carry[9] , \add_66/carry[8] , \add_66/carry[7] ,
         \add_66/carry[6] , \add_66/carry[5] , \add_66/carry[4] ,
         \add_66/carry[3] , \add_66/carry[2] , n3, n13, n15, n16, n17, n18,
         n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n261, n263, n264, n265, n266, n267, n269, n270, n272, n273, n274,
         n275, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292;
  assign \U11/DATA1_0  = ReadBus[0];
  assign \U11/DATA1_1  = ReadBus[1];
  assign \U11/DATA1_2  = ReadBus[2];
  assign \U11/DATA1_3  = ReadBus[3];
  assign \U11/DATA1_4  = ReadBus[4];
  assign \U11/DATA1_5  = ReadBus[5];
  assign \U11/DATA1_6  = ReadBus[6];
  assign \U11/DATA1_7  = ReadBus[7];
  assign \U11/DATA1_8  = ReadBus[8];
  assign \U11/DATA1_9  = ReadBus[9];
  assign \U11/DATA1_10  = ReadBus[10];
  assign \U11/DATA1_11  = ReadBus[11];
  assign \U11/DATA1_12  = ReadBus[12];
  assign \U11/DATA1_13  = ReadBus[13];
  assign \U11/DATA1_14  = ReadBus[14];
  assign \U11/DATA1_15  = ReadBus[15];
  assign \U11/DATA1_16  = ReadBus[16];
  assign \U11/DATA1_17  = ReadBus[17];
  assign \U11/DATA1_18  = ReadBus[18];
  assign \U11/DATA1_19  = ReadBus[19];
  assign ReadAddr[0] = \U10/DATA1_0 ;
  assign ReadAddr[1] = \U10/DATA1_1 ;
  assign ReadAddr[2] = \U10/DATA1_2 ;
  assign ReadAddr[3] = \U10/DATA1_3 ;
  assign ReadAddr[4] = \U10/DATA1_4 ;
  assign ReadAddr[5] = \U10/DATA1_5 ;
  assign ReadAddr[6] = \U10/DATA1_6 ;
  assign ReadAddr[7] = \U10/DATA1_7 ;
  assign ReadAddr[8] = \U10/DATA1_8 ;
  assign ReadAddr[9] = \U10/DATA1_9 ;
  assign ReadAddr[10] = \U10/DATA1_10 ;
  assign ReadAddr[11] = \U10/DATA1_11 ;
  assign ReadAddr[12] = \U10/DATA1_12 ;
  assign ReadAddr[13] = \U10/DATA1_13 ;
  assign ReadAddr[14] = \U10/DATA1_14 ;
  assign ReadAddr[15] = \U10/DATA1_15 ;
  assign \U4/DATA3_0  = input_base_offset;

  HA_X1 \add_66/U1_1_1  ( .A(\U10/DATA1_1 ), .B(\U10/DATA1_0 ), .CO(
        \add_66/carry[2] ), .S(\U5/DATA1_1 ) );
  HA_X1 \add_66/U1_1_2  ( .A(\U10/DATA1_2 ), .B(\add_66/carry[2] ), .CO(
        \add_66/carry[3] ), .S(\U5/DATA1_2 ) );
  HA_X1 \add_66/U1_1_3  ( .A(\U10/DATA1_3 ), .B(\add_66/carry[3] ), .CO(
        \add_66/carry[4] ), .S(\U5/DATA1_3 ) );
  HA_X1 \add_66/U1_1_4  ( .A(\U10/DATA1_4 ), .B(\add_66/carry[4] ), .CO(
        \add_66/carry[5] ), .S(\U5/DATA1_4 ) );
  HA_X1 \add_66/U1_1_5  ( .A(\U10/DATA1_5 ), .B(\add_66/carry[5] ), .CO(
        \add_66/carry[6] ), .S(\U5/DATA1_5 ) );
  HA_X1 \add_66/U1_1_6  ( .A(\U10/DATA1_6 ), .B(\add_66/carry[6] ), .CO(
        \add_66/carry[7] ), .S(\U5/DATA1_6 ) );
  HA_X1 \add_66/U1_1_7  ( .A(\U10/DATA1_7 ), .B(\add_66/carry[7] ), .CO(
        \add_66/carry[8] ), .S(\U5/DATA1_7 ) );
  HA_X1 \add_66/U1_1_8  ( .A(\U10/DATA1_8 ), .B(\add_66/carry[8] ), .CO(
        \add_66/carry[9] ), .S(\U5/DATA1_8 ) );
  HA_X1 \add_66/U1_1_9  ( .A(\U10/DATA1_9 ), .B(\add_66/carry[9] ), .CO(
        \add_66/carry[10] ), .S(\U5/DATA1_9 ) );
  HA_X1 \add_66/U1_1_10  ( .A(\U10/DATA1_10 ), .B(\add_66/carry[10] ), .CO(
        \add_66/carry[11] ), .S(\U5/DATA1_10 ) );
  HA_X1 \add_66/U1_1_11  ( .A(\U10/DATA1_11 ), .B(\add_66/carry[11] ), .CO(
        \add_66/carry[12] ), .S(\U5/DATA1_11 ) );
  HA_X1 \add_66/U1_1_13  ( .A(n261), .B(\U10/DATA1_13 ), .CO(
        \add_66/carry[14] ), .S(\U5/DATA1_13 ) );
  HA_X1 \add_69/U1_1_1  ( .A(\add_69/A[1] ), .B(\add_69/A[0] ), .CO(
        \add_69/carry[2] ), .S(\U3/U1/DATA1_1 ) );
  HA_X1 \add_69/U1_1_2  ( .A(\add_69/A[2] ), .B(\add_69/carry[2] ), .CO(
        \add_69/carry[3] ), .S(\U3/U1/DATA1_2 ) );
  HA_X1 \add_69/U1_1_3  ( .A(\add_69/A[3] ), .B(\add_69/carry[3] ), .CO(
        \add_69/carry[4] ), .S(\U3/U1/DATA1_3 ) );
  HA_X1 \add_69/U1_1_4  ( .A(\add_69/A[4] ), .B(\add_69/carry[4] ), .CO(
        \add_69/carry[5] ), .S(\U3/U1/DATA1_4 ) );
  HA_X1 \add_69/U1_1_5  ( .A(\add_69/A[5] ), .B(\add_69/carry[5] ), .CO(
        \add_69/carry[6] ), .S(\U3/U1/DATA1_5 ) );
  HA_X1 \add_69/U1_1_6  ( .A(\add_69/A[6] ), .B(\add_69/carry[6] ), .CO(
        \add_69/carry[7] ), .S(\U3/U1/DATA1_6 ) );
  HA_X1 \add_69/U1_1_7  ( .A(\add_69/A[7] ), .B(\add_69/carry[7] ), .CO(
        \add_69/carry[8] ), .S(\U3/U1/DATA1_7 ) );
  DFFR_X1 \count_reg[0]  ( .D(n33), .CK(clock), .RN(n281), .Q(\add_69/A[0] ), 
        .QN(n13) );
  DFFR_X1 \count_reg[8]  ( .D(n32), .CK(clock), .RN(n279), .Q(\add_69/A[8] ), 
        .QN(n3) );
  DFFR_X1 \ReadAddress_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .RN(n279), .Q(
        \U10/DATA1_1 ) );
  DFFR_X1 \StoreAddress_reg[1]  ( .D(\U10/Z_1 ), .CK(clock), .RN(n279), .Q(
        StoreAddress[1]) );
  DFFR_X1 \ReadAddress_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .RN(n279), .Q(
        \U10/DATA1_2 ) );
  DFFR_X1 \StoreAddress_reg[2]  ( .D(\U10/Z_2 ), .CK(clock), .RN(n279), .Q(
        StoreAddress[2]) );
  DFFR_X1 \ReadAddress_reg[3]  ( .D(\U5/Z_3 ), .CK(clock), .RN(n279), .Q(
        \U10/DATA1_3 ) );
  DFFR_X1 \StoreAddress_reg[3]  ( .D(\U10/Z_3 ), .CK(clock), .RN(n279), .Q(
        StoreAddress[3]) );
  DFFR_X1 \ReadAddress_reg[4]  ( .D(\U5/Z_4 ), .CK(clock), .RN(n279), .Q(
        \U10/DATA1_4 ) );
  DFFR_X1 \StoreAddress_reg[4]  ( .D(\U10/Z_4 ), .CK(clock), .RN(n279), .Q(
        StoreAddress[4]) );
  DFFR_X1 \ReadAddress_reg[5]  ( .D(\U5/Z_5 ), .CK(clock), .RN(n279), .Q(
        \U10/DATA1_5 ) );
  DFFR_X1 \StoreAddress_reg[5]  ( .D(\U10/Z_5 ), .CK(clock), .RN(n280), .Q(
        StoreAddress[5]) );
  DFFR_X1 \ReadAddress_reg[6]  ( .D(\U5/Z_6 ), .CK(clock), .RN(n280), .Q(
        \U10/DATA1_6 ) );
  DFFR_X1 \StoreAddress_reg[6]  ( .D(\U10/Z_6 ), .CK(clock), .RN(n280), .Q(
        StoreAddress[6]) );
  DFFR_X1 \ReadAddress_reg[7]  ( .D(\U5/Z_7 ), .CK(clock), .RN(n280), .Q(
        \U10/DATA1_7 ) );
  DFFR_X1 \StoreAddress_reg[7]  ( .D(\U10/Z_7 ), .CK(clock), .RN(n280), .Q(
        StoreAddress[7]) );
  DFFR_X1 \ReadAddress_reg[8]  ( .D(\U5/Z_8 ), .CK(clock), .RN(n280), .Q(
        \U10/DATA1_8 ) );
  DFFR_X1 \StoreAddress_reg[8]  ( .D(\U10/Z_8 ), .CK(clock), .RN(n280), .Q(
        StoreAddress[8]) );
  DFFR_X1 \ReadAddress_reg[9]  ( .D(\U5/Z_9 ), .CK(clock), .RN(n280), .Q(
        \U10/DATA1_9 ) );
  DFFR_X1 \StoreAddress_reg[9]  ( .D(\U10/Z_9 ), .CK(clock), .RN(n280), .Q(
        StoreAddress[9]) );
  DFFR_X1 \ReadAddress_reg[10]  ( .D(\U5/Z_10 ), .CK(clock), .RN(n280), .Q(
        \U10/DATA1_10 ) );
  DFFR_X1 \StoreAddress_reg[10]  ( .D(\U10/Z_10 ), .CK(clock), .RN(n280), .Q(
        StoreAddress[10]) );
  DFFR_X1 \ReadAddress_reg[11]  ( .D(\U5/Z_11 ), .CK(clock), .RN(n280), .Q(
        \U10/DATA1_11 ) );
  DFFR_X1 \StoreAddress_reg[11]  ( .D(\U10/Z_11 ), .CK(clock), .RN(n281), .Q(
        StoreAddress[11]) );
  DFFR_X1 \ReadAddress_reg[12]  ( .D(\U5/Z_12 ), .CK(clock), .RN(n281), .Q(
        \U10/DATA1_12 ) );
  DFFR_X1 \StoreAddress_reg[12]  ( .D(\U10/Z_12 ), .CK(clock), .RN(n281), .Q(
        StoreAddress[12]) );
  DFFR_X1 \ReadAddress_reg[13]  ( .D(\U5/Z_13 ), .CK(clock), .RN(n281), .Q(
        \U10/DATA1_13 ) );
  DFFR_X1 \StoreAddress_reg[13]  ( .D(\U10/Z_13 ), .CK(clock), .RN(n281), .Q(
        StoreAddress[13]) );
  DFFR_X1 \StoreAddress_reg[14]  ( .D(\U10/Z_14 ), .CK(clock), .RN(n281), .Q(
        StoreAddress[14]) );
  DFFR_X1 \StoreAddress_reg[0]  ( .D(\U10/Z_0 ), .CK(clock), .RN(n281), .Q(
        StoreAddress[0]) );
  DFFR_X1 \StoreAddress_reg[15]  ( .D(\U10/Z_15 ), .CK(clock), .RN(n281), .Q(
        StoreAddress[15]) );
  DFFR_X1 \count_reg[1]  ( .D(n291), .CK(clock), .RN(n281), .Q(\add_69/A[1] )
         );
  DFFR_X1 \count_reg[2]  ( .D(n290), .CK(clock), .RN(n282), .Q(\add_69/A[2] )
         );
  DFFR_X1 \count_reg[3]  ( .D(n289), .CK(clock), .RN(n282), .Q(\add_69/A[3] )
         );
  DFFR_X1 \count_reg[4]  ( .D(n288), .CK(clock), .RN(n282), .Q(\add_69/A[4] )
         );
  DFFR_X1 \count_reg[5]  ( .D(n287), .CK(clock), .RN(n282), .Q(\add_69/A[5] )
         );
  DFFR_X1 \count_reg[6]  ( .D(n286), .CK(clock), .RN(n282), .Q(\add_69/A[6] )
         );
  DFFR_X1 \count_reg[7]  ( .D(n285), .CK(clock), .RN(n282), .Q(\add_69/A[7] )
         );
  SDFFR_X2 StartOut_reg ( .D(1'b0), .SI(start), .SE(n3), .CK(clock), .RN(
        reset_n), .Q(StartOut) );
  DFFR_X1 \AccumlateOut_reg[19]  ( .D(\U7/Z_19 ), .CK(clock), .RN(n282), .Q(
        AccumlateOut[19]) );
  DFFR_X1 \AccumlateOut_reg[18]  ( .D(\U7/Z_18 ), .CK(clock), .RN(n282), .Q(
        AccumlateOut[18]) );
  DFFR_X1 \AccumlateOut_reg[17]  ( .D(\U7/Z_17 ), .CK(clock), .RN(n282), .Q(
        AccumlateOut[17]) );
  DFFR_X1 \AccumlateOut_reg[16]  ( .D(\U7/Z_16 ), .CK(clock), .RN(n282), .Q(
        AccumlateOut[16]) );
  DFFR_X1 \AccumlateOut_reg[15]  ( .D(\U7/Z_15 ), .CK(clock), .RN(n282), .Q(
        AccumlateOut[15]) );
  DFFR_X1 \AccumlateOut_reg[14]  ( .D(\U7/Z_14 ), .CK(clock), .RN(n282), .Q(
        AccumlateOut[14]) );
  DFFR_X1 \AccumlateOut_reg[13]  ( .D(\U7/Z_13 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[13]) );
  DFFR_X1 \AccumlateOut_reg[12]  ( .D(\U7/Z_12 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[12]) );
  DFFR_X1 \AccumlateOut_reg[11]  ( .D(\U7/Z_11 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[11]) );
  DFFR_X1 \AccumlateOut_reg[10]  ( .D(\U7/Z_10 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[10]) );
  DFFR_X1 \AccumlateOut_reg[9]  ( .D(\U7/Z_9 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[9]) );
  DFFR_X1 \AccumlateOut_reg[8]  ( .D(\U7/Z_8 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[8]) );
  DFFR_X1 \AccumlateOut_reg[7]  ( .D(\U7/Z_7 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[7]) );
  DFFR_X1 \AccumlateOut_reg[6]  ( .D(\U7/Z_6 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[6]) );
  DFFR_X1 \AccumlateOut_reg[5]  ( .D(\U7/Z_5 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[5]) );
  DFFR_X1 \AccumlateOut_reg[0]  ( .D(\U7/Z_0 ), .CK(clock), .RN(reset_n), .Q(
        AccumlateOut[0]) );
  SDFFR_X2 done0_reg ( .D(1'b0), .SI(\add_69/A[8] ), .SE(start), .CK(clock), 
        .RN(reset_n), .Q(\U9/DATA1_0 ) );
  DFFR_X1 done1_reg ( .D(\U9/Z_0 ), .CK(clock), .RN(reset_n), .Q(\U8/DATA1_0 )
         );
  DFFR_X1 done_reg ( .D(\U8/Z_0 ), .CK(clock), .RN(n279), .Q(done) );
  NAND2_X2 U12 ( .A1(n292), .A2(n22), .ZN(n32) );
  NAND2_X2 U13 ( .A1(\add_69/carry[8] ), .A2(n277), .ZN(n22) );
  OAI22_X2 U14 ( .A1(n292), .A2(n13), .B1(\add_69/A[0] ), .B2(n264), .ZN(n33)
         );
  NOR2_X2 U16 ( .A1(n28), .A2(n29), .ZN(n27) );
  NAND4_X2 U17 ( .A1(ReadBus[35]), .A2(ReadBus[33]), .A3(ReadBus[31]), .A4(
        ReadBus[29]), .ZN(n29) );
  NAND4_X2 U18 ( .A1(ReadBus[27]), .A2(ReadBus[25]), .A3(ReadBus[23]), .A4(
        ReadBus[21]), .ZN(n28) );
  NOR4_X2 U19 ( .A1(ReadBus[24]), .A2(ReadBus[22]), .A3(ReadBus[20]), .A4(n278), .ZN(n26) );
  NOR3_X2 U20 ( .A1(ReadBus[30]), .A2(ReadBus[34]), .A3(ReadBus[32]), .ZN(n25)
         );
  NOR2_X2 U21 ( .A1(ReadBus[28]), .A2(ReadBus[26]), .ZN(n24) );
  NAND2_X2 U24 ( .A1(\U4/DATA3_0 ), .A2(n278), .ZN(n31) );
  NOR2_X2 U26 ( .A1(n278), .A2(n277), .ZN(\U4/CONTROL2 ) );
  AND2_X1 U38 ( .A1(\U9/DATA1_0 ), .A2(start), .ZN(\U9/Z_0 ) );
  AND2_X1 U39 ( .A1(\U8/DATA1_0 ), .A2(start), .ZN(\U8/Z_0 ) );
  AND2_X1 U48 ( .A1(\U11/DATA1_19 ), .A2(n263), .ZN(\U7/Z_19 ) );
  AND2_X1 U49 ( .A1(\U11/DATA1_18 ), .A2(n263), .ZN(\U7/Z_18 ) );
  AND2_X1 U50 ( .A1(\U11/DATA1_17 ), .A2(n263), .ZN(\U7/Z_17 ) );
  AND2_X1 U51 ( .A1(\U11/DATA1_16 ), .A2(n263), .ZN(\U7/Z_16 ) );
  AND2_X1 U52 ( .A1(\U11/DATA1_15 ), .A2(n263), .ZN(\U7/Z_15 ) );
  AND2_X1 U53 ( .A1(\U11/DATA1_14 ), .A2(n263), .ZN(\U7/Z_14 ) );
  AND2_X1 U54 ( .A1(\U11/DATA1_13 ), .A2(n263), .ZN(\U7/Z_13 ) );
  AND2_X1 U60 ( .A1(\U5/DATA1_9 ), .A2(n277), .ZN(\U5/Z_9 ) );
  AND2_X1 U61 ( .A1(\U5/DATA1_8 ), .A2(n277), .ZN(\U5/Z_8 ) );
  AND2_X1 U62 ( .A1(\U5/DATA1_7 ), .A2(n277), .ZN(\U5/Z_7 ) );
  AND2_X1 U63 ( .A1(\U5/DATA1_6 ), .A2(n277), .ZN(\U5/Z_6 ) );
  AND2_X1 U64 ( .A1(\U5/DATA1_5 ), .A2(n277), .ZN(\U5/Z_5 ) );
  AND2_X1 U65 ( .A1(\U5/DATA1_4 ), .A2(n277), .ZN(\U5/Z_4 ) );
  AND2_X1 U66 ( .A1(\U5/DATA1_3 ), .A2(n277), .ZN(\U5/Z_3 ) );
  AND2_X1 U67 ( .A1(\U5/DATA1_2 ), .A2(n277), .ZN(\U5/Z_2 ) );
  AND2_X1 U68 ( .A1(\U5/DATA1_14 ), .A2(n277), .ZN(\U5/Z_14 ) );
  AND2_X1 U69 ( .A1(\U5/DATA1_13 ), .A2(n277), .ZN(\U5/Z_13 ) );
  AND2_X1 U70 ( .A1(\U5/DATA1_12 ), .A2(n277), .ZN(\U5/Z_12 ) );
  AND2_X1 U71 ( .A1(\U5/DATA1_11 ), .A2(n277), .ZN(\U5/Z_11 ) );
  AND2_X1 U72 ( .A1(\U5/DATA1_10 ), .A2(n277), .ZN(\U5/Z_10 ) );
  AND2_X1 U73 ( .A1(\U5/DATA1_1 ), .A2(n277), .ZN(\U5/Z_1 ) );
  AND2_X1 U74 ( .A1(\U10/DATA1_9 ), .A2(start), .ZN(\U10/Z_9 ) );
  AND2_X1 U75 ( .A1(\U10/DATA1_8 ), .A2(start), .ZN(\U10/Z_8 ) );
  AND2_X1 U76 ( .A1(\U10/DATA1_7 ), .A2(start), .ZN(\U10/Z_7 ) );
  AND2_X1 U77 ( .A1(\U10/DATA1_6 ), .A2(start), .ZN(\U10/Z_6 ) );
  AND2_X1 U78 ( .A1(\U10/DATA1_5 ), .A2(start), .ZN(\U10/Z_5 ) );
  AND2_X1 U79 ( .A1(\U10/DATA1_4 ), .A2(start), .ZN(\U10/Z_4 ) );
  AND2_X1 U80 ( .A1(\U10/DATA1_3 ), .A2(start), .ZN(\U10/Z_3 ) );
  AND2_X1 U81 ( .A1(\U10/DATA1_2 ), .A2(start), .ZN(\U10/Z_2 ) );
  AND2_X1 U82 ( .A1(start), .A2(\U10/DATA1_15 ), .ZN(\U10/Z_15 ) );
  AND2_X1 U83 ( .A1(\U10/DATA1_14 ), .A2(start), .ZN(\U10/Z_14 ) );
  AND2_X1 U84 ( .A1(\U10/DATA1_13 ), .A2(start), .ZN(\U10/Z_13 ) );
  AND2_X1 U85 ( .A1(\U10/DATA1_12 ), .A2(start), .ZN(\U10/Z_12 ) );
  AND2_X1 U86 ( .A1(\U10/DATA1_11 ), .A2(start), .ZN(\U10/Z_11 ) );
  AND2_X1 U87 ( .A1(\U10/DATA1_10 ), .A2(start), .ZN(\U10/Z_10 ) );
  AND2_X1 U88 ( .A1(\U10/DATA1_1 ), .A2(start), .ZN(\U10/Z_1 ) );
  AND2_X1 U89 ( .A1(start), .A2(\U10/DATA1_0 ), .ZN(\U10/Z_0 ) );
  DFFR_X2 \AccumlateOut_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .RN(n283), .QN(
        n267) );
  DFFR_X2 \AccumlateOut_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .RN(reset_n), .QN(
        n270) );
  DFFR_X2 \ReadAddress_reg[14]  ( .D(\U5/Z_14 ), .CK(clock), .RN(n281), .Q(
        \U10/DATA1_14 ), .QN(n266) );
  DFFR_X2 \AccumlateOut_reg[4]  ( .D(\U7/Z_4 ), .CK(clock), .RN(n283), .Q(
        AccumlateOut[4]) );
  DFFR_X2 \AccumlateOut_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .RN(reset_n), .QN(
        n275) );
  DFFR_X2 \ReadAddress_reg[0]  ( .D(\U5/Z_0 ), .CK(clock), .RN(n279), .Q(
        \U10/DATA1_0 ) );
  DFFR_X2 \ReadAddress_reg[15]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n281), .Q(
        \U10/DATA1_15 ), .QN(n272) );
  AND2_X4 U5 ( .A1(\U10/DATA1_12 ), .A2(\add_66/carry[12] ), .ZN(n261) );
  AND4_X4 U6 ( .A1(n26), .A2(n27), .A3(n24), .A4(n25), .ZN(n263) );
  OR2_X4 U7 ( .A1(\add_69/A[8] ), .A2(n278), .ZN(n264) );
  XOR2_X2 U8 ( .A(\U10/DATA1_12 ), .B(\add_66/carry[12] ), .Z(\U5/DATA1_12 )
         );
  AND2_X1 U9 ( .A1(\U10/DATA1_13 ), .A2(n261), .ZN(n265) );
  NAND2_X2 U10 ( .A1(\U10/DATA1_14 ), .A2(n265), .ZN(n269) );
  XNOR2_X1 U11 ( .A(n266), .B(\add_66/carry[14] ), .ZN(\U5/DATA1_14 ) );
  INV_X4 U15 ( .A(n267), .ZN(AccumlateOut[2]) );
  INV_X2 U22 ( .A(n269), .ZN(\add_66/carry[15] ) );
  NAND2_X2 U23 ( .A1(\U10/DATA1_15 ), .A2(\add_66/carry[15] ), .ZN(n273) );
  INV_X4 U25 ( .A(n270), .ZN(AccumlateOut[3]) );
  NAND2_X2 U27 ( .A1(n272), .A2(n269), .ZN(n274) );
  NAND2_X2 U28 ( .A1(n273), .A2(n274), .ZN(n30) );
  INV_X4 U29 ( .A(n275), .ZN(AccumlateOut[1]) );
  NOR2_X1 U30 ( .A1(\U10/DATA1_0 ), .A2(n264), .ZN(\U5/Z_0 ) );
  INV_X4 U31 ( .A(n284), .ZN(n282) );
  INV_X4 U32 ( .A(n284), .ZN(n280) );
  INV_X4 U33 ( .A(n284), .ZN(n279) );
  INV_X4 U34 ( .A(n284), .ZN(n281) );
  INV_X4 U35 ( .A(n284), .ZN(n283) );
  INV_X4 U36 ( .A(start), .ZN(n278) );
  INV_X4 U37 ( .A(reset_n), .ZN(n284) );
  INV_X4 U40 ( .A(n264), .ZN(n277) );
  OAI21_X2 U41 ( .B1(n30), .B2(n264), .A(n31), .ZN(\U4/Z_0 ) );
  AOI22_X2 U42 ( .A1(\U3/U1/DATA1_7 ), .A2(n277), .B1(\add_69/A[7] ), .B2(
        \U4/CONTROL2 ), .ZN(n21) );
  AOI22_X2 U43 ( .A1(\U3/U1/DATA1_6 ), .A2(n277), .B1(\add_69/A[6] ), .B2(
        \U4/CONTROL2 ), .ZN(n20) );
  AOI22_X2 U44 ( .A1(\U3/U1/DATA1_5 ), .A2(n277), .B1(\add_69/A[5] ), .B2(
        \U4/CONTROL2 ), .ZN(n19) );
  AOI22_X2 U45 ( .A1(\U3/U1/DATA1_4 ), .A2(n277), .B1(\add_69/A[4] ), .B2(
        \U4/CONTROL2 ), .ZN(n18) );
  AOI22_X2 U46 ( .A1(\U3/U1/DATA1_3 ), .A2(n277), .B1(\add_69/A[3] ), .B2(
        \U4/CONTROL2 ), .ZN(n17) );
  AOI22_X2 U47 ( .A1(\U3/U1/DATA1_2 ), .A2(n277), .B1(\add_69/A[2] ), .B2(
        \U4/CONTROL2 ), .ZN(n16) );
  AOI22_X2 U55 ( .A1(\U3/U1/DATA1_1 ), .A2(n277), .B1(\add_69/A[1] ), .B2(
        \U4/CONTROL2 ), .ZN(n15) );
  AND2_X1 U56 ( .A1(\U11/DATA1_0 ), .A2(n263), .ZN(\U7/Z_0 ) );
  AND2_X1 U57 ( .A1(\U11/DATA1_1 ), .A2(n263), .ZN(\U7/Z_1 ) );
  AND2_X1 U58 ( .A1(\U11/DATA1_2 ), .A2(n263), .ZN(\U7/Z_2 ) );
  AND2_X1 U59 ( .A1(\U11/DATA1_3 ), .A2(n263), .ZN(\U7/Z_3 ) );
  AND2_X1 U90 ( .A1(\U11/DATA1_4 ), .A2(n263), .ZN(\U7/Z_4 ) );
  AND2_X1 U91 ( .A1(\U11/DATA1_5 ), .A2(n263), .ZN(\U7/Z_5 ) );
  AND2_X1 U92 ( .A1(\U11/DATA1_6 ), .A2(n263), .ZN(\U7/Z_6 ) );
  AND2_X1 U93 ( .A1(\U11/DATA1_7 ), .A2(n263), .ZN(\U7/Z_7 ) );
  AND2_X1 U94 ( .A1(\U11/DATA1_8 ), .A2(n263), .ZN(\U7/Z_8 ) );
  AND2_X1 U95 ( .A1(\U11/DATA1_9 ), .A2(n263), .ZN(\U7/Z_9 ) );
  AND2_X1 U96 ( .A1(\U11/DATA1_10 ), .A2(n263), .ZN(\U7/Z_10 ) );
  AND2_X1 U97 ( .A1(\U11/DATA1_11 ), .A2(n263), .ZN(\U7/Z_11 ) );
  AND2_X1 U98 ( .A1(\U11/DATA1_12 ), .A2(n263), .ZN(\U7/Z_12 ) );
  INV_X4 U99 ( .A(n21), .ZN(n285) );
  INV_X4 U100 ( .A(n20), .ZN(n286) );
  INV_X4 U101 ( .A(n19), .ZN(n287) );
  INV_X4 U102 ( .A(n18), .ZN(n288) );
  INV_X4 U103 ( .A(n17), .ZN(n289) );
  INV_X4 U104 ( .A(n16), .ZN(n290) );
  INV_X4 U105 ( .A(n15), .ZN(n291) );
  INV_X4 U106 ( .A(\U4/CONTROL2 ), .ZN(n292) );
endmodule


module Cdf_Accumlate ( clock, reset_n, AccumlateIn, StartIn, StoreAddressIn, 
        AccumlateResult, StoreAddressOut, StartOut, CdfMin, CdfValid );
  input [19:0] AccumlateIn;
  input [15:0] StoreAddressIn;
  output [19:0] AccumlateResult;
  output [15:0] StoreAddressOut;
  output [19:0] CdfMin;
  input clock, reset_n, StartIn;
  output StartOut, CdfValid;
  wire   \U8/Z_0 , \U6/DATA2_0 , \U6/DATA2_1 , \U6/DATA2_2 , \U6/DATA2_3 ,
         \U6/DATA2_4 , \U6/DATA2_5 , \U6/DATA2_6 , \U6/DATA2_7 , \U6/DATA2_8 ,
         \U6/DATA2_9 , \U6/DATA2_10 , \U6/DATA2_11 , \U6/DATA2_12 ,
         \U6/DATA2_13 , \U6/DATA2_14 , \U6/DATA2_15 , \U6/DATA2_16 ,
         \U6/DATA2_17 , \U6/DATA2_18 , \U6/DATA2_19 , \U6/DATA1_2 ,
         \U6/DATA1_3 , \U6/DATA1_4 , \U6/DATA1_5 , \U6/DATA1_6 , \U6/DATA1_7 ,
         \U6/DATA1_10 , \U6/DATA1_11 , \U6/DATA1_12 , \U6/DATA1_13 ,
         \U6/DATA1_14 , \U6/DATA1_15 , \add/B[0] , \add/B[1] , \add/B[2] ,
         \add/B[3] , \add/B[4] , \add/B[5] , \add/B[6] , \add/B[7] ,
         \add/B[8] , \add/B[9] , \add/B[10] , \add/B[11] , \add/B[12] ,
         \add/B[13] , \add/B[14] , \add/B[15] , \add/B[16] , \add/B[17] ,
         \add/B[18] , \add/B[19] , \add/A[0] , \add/A[1] , \add/A[2] ,
         \add/A[3] , \add/A[4] , \add/A[5] , \add/A[6] , \add/A[7] ,
         \add/A[8] , \add/A[9] , \add/A[10] , \add/A[11] , \add/A[12] ,
         \add/A[13] , \add/A[14] , \add/A[15] , \add/A[16] , \add/A[17] ,
         \add/A[18] , \add/A[19] , n76, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n242, n243, n244,
         n245, n246, n247, n248, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454;
  assign CdfMin[0] = \U6/DATA2_0 ;
  assign CdfMin[1] = \U6/DATA2_1 ;
  assign CdfMin[2] = \U6/DATA2_2 ;
  assign CdfMin[3] = \U6/DATA2_3 ;
  assign CdfMin[4] = \U6/DATA2_4 ;
  assign CdfMin[5] = \U6/DATA2_5 ;
  assign CdfMin[6] = \U6/DATA2_6 ;
  assign CdfMin[7] = \U6/DATA2_7 ;
  assign CdfMin[8] = \U6/DATA2_8 ;
  assign CdfMin[9] = \U6/DATA2_9 ;
  assign CdfMin[10] = \U6/DATA2_10 ;
  assign CdfMin[11] = \U6/DATA2_11 ;
  assign CdfMin[12] = \U6/DATA2_12 ;
  assign CdfMin[13] = \U6/DATA2_13 ;
  assign CdfMin[14] = \U6/DATA2_14 ;
  assign CdfMin[15] = \U6/DATA2_15 ;
  assign CdfMin[16] = \U6/DATA2_16 ;
  assign CdfMin[17] = \U6/DATA2_17 ;
  assign CdfMin[18] = \U6/DATA2_18 ;
  assign CdfMin[19] = \U6/DATA2_19 ;
  assign \add/B[0]  = AccumlateIn[0];
  assign \add/B[1]  = AccumlateIn[1];
  assign \add/B[2]  = AccumlateIn[2];
  assign \add/B[3]  = AccumlateIn[3];
  assign \add/B[4]  = AccumlateIn[4];
  assign \add/B[5]  = AccumlateIn[5];
  assign \add/B[6]  = AccumlateIn[6];
  assign \add/B[7]  = AccumlateIn[7];
  assign \add/B[8]  = AccumlateIn[8];
  assign \add/B[9]  = AccumlateIn[9];
  assign \add/B[10]  = AccumlateIn[10];
  assign \add/B[11]  = AccumlateIn[11];
  assign \add/B[12]  = AccumlateIn[12];
  assign \add/B[13]  = AccumlateIn[13];
  assign \add/B[14]  = AccumlateIn[14];
  assign \add/B[15]  = AccumlateIn[15];
  assign \add/B[16]  = AccumlateIn[16];
  assign \add/B[17]  = AccumlateIn[17];
  assign \add/B[18]  = AccumlateIn[18];
  assign \add/B[19]  = AccumlateIn[19];
  assign AccumlateResult[0] = \add/A[0] ;
  assign AccumlateResult[1] = \add/A[1] ;
  assign AccumlateResult[2] = \add/A[2] ;
  assign AccumlateResult[3] = \add/A[3] ;
  assign AccumlateResult[4] = \add/A[4] ;
  assign AccumlateResult[5] = \add/A[5] ;
  assign AccumlateResult[6] = \add/A[6] ;
  assign AccumlateResult[7] = \add/A[7] ;
  assign AccumlateResult[8] = \add/A[8] ;
  assign AccumlateResult[9] = \add/A[9] ;
  assign AccumlateResult[10] = \add/A[10] ;
  assign AccumlateResult[11] = \add/A[11] ;
  assign AccumlateResult[12] = \add/A[12] ;
  assign AccumlateResult[13] = \add/A[13] ;
  assign AccumlateResult[14] = \add/A[14] ;
  assign AccumlateResult[15] = \add/A[15] ;
  assign AccumlateResult[16] = \add/A[16] ;
  assign AccumlateResult[17] = \add/A[17] ;
  assign AccumlateResult[18] = \add/A[18] ;
  assign AccumlateResult[19] = \add/A[19] ;

  DFFR_X1 \AccumlateResult_reg[0]  ( .D(n240), .CK(clock), .RN(n310), .Q(
        \add/A[0] ), .QN(n253) );
  SDFFR_X2 \AccumlateResult_reg[2]  ( .D(1'b0), .SI(StartIn), .SE(\U6/DATA1_2 ), .CK(clock), .RN(reset_n), .Q(\add/A[2] ), .QN(n220) );
  SDFFR_X2 \AccumlateResult_reg[3]  ( .D(1'b0), .SI(StartIn), .SE(\U6/DATA1_3 ), .CK(clock), .RN(reset_n), .Q(\add/A[3] ) );
  SDFFR_X2 \AccumlateResult_reg[4]  ( .D(1'b0), .SI(StartIn), .SE(\U6/DATA1_4 ), .CK(clock), .RN(reset_n), .Q(\add/A[4] ) );
  SDFFR_X2 \AccumlateResult_reg[6]  ( .D(1'b0), .SI(StartIn), .SE(\U6/DATA1_6 ), .CK(clock), .RN(reset_n), .Q(\add/A[6] ) );
  SDFFR_X2 \AccumlateResult_reg[7]  ( .D(1'b0), .SI(StartIn), .SE(\U6/DATA1_7 ), .CK(clock), .RN(reset_n), .Q(\add/A[7] ) );
  DFFR_X1 \AccumlateResult_reg[8]  ( .D(n232), .CK(clock), .RN(n310), .Q(
        \add/A[8] ) );
  SDFFR_X2 \AccumlateResult_reg[10]  ( .D(1'b0), .SI(StartIn), .SE(
        \U6/DATA1_10 ), .CK(clock), .RN(reset_n), .Q(\add/A[10] ), .QN(n223)
         );
  SDFFR_X2 \AccumlateResult_reg[11]  ( .D(1'b0), .SI(StartIn), .SE(
        \U6/DATA1_11 ), .CK(clock), .RN(reset_n), .Q(\add/A[11] ), .QN(n222)
         );
  SDFFR_X2 \AccumlateResult_reg[12]  ( .D(1'b0), .SI(StartIn), .SE(
        \U6/DATA1_12 ), .CK(clock), .RN(reset_n), .Q(\add/A[12] ), .QN(n224)
         );
  SDFFR_X2 \AccumlateResult_reg[13]  ( .D(1'b0), .SI(StartIn), .SE(
        \U6/DATA1_13 ), .CK(clock), .RN(reset_n), .Q(\add/A[13] ), .QN(n221)
         );
  SDFFR_X2 \AccumlateResult_reg[14]  ( .D(1'b0), .SI(StartIn), .SE(
        \U6/DATA1_14 ), .CK(clock), .RN(reset_n), .Q(\add/A[14] ), .QN(n227)
         );
  SDFFR_X2 \AccumlateResult_reg[15]  ( .D(1'b0), .SI(StartIn), .SE(
        \U6/DATA1_15 ), .CK(clock), .RN(reset_n), .Q(\add/A[15] ), .QN(n225)
         );
  DFFR_X1 \AccumlateResult_reg[16]  ( .D(n287), .CK(clock), .RN(n310), .Q(
        \add/A[16] ), .QN(n234) );
  DFFR_X1 \AccumlateResult_reg[17]  ( .D(n286), .CK(clock), .RN(n310), .Q(
        \add/A[17] ) );
  DFFR_X1 \AccumlateResult_reg[18]  ( .D(n302), .CK(clock), .RN(n310), .Q(
        \add/A[18] ), .QN(n236) );
  DFFR_X1 \CdfMin_reg[0]  ( .D(n454), .CK(clock), .RN(n310), .Q(\U6/DATA2_0 ), 
        .QN(n229) );
  DFFR_X1 \CdfMin_reg[1]  ( .D(n453), .CK(clock), .RN(n310), .Q(\U6/DATA2_1 ), 
        .QN(n238) );
  DFFR_X1 \CdfMin_reg[2]  ( .D(n452), .CK(clock), .RN(n311), .Q(\U6/DATA2_2 ), 
        .QN(n248) );
  DFFR_X1 \CdfMin_reg[3]  ( .D(n451), .CK(clock), .RN(n311), .Q(\U6/DATA2_3 ), 
        .QN(n246) );
  DFFR_X1 \CdfMin_reg[4]  ( .D(n450), .CK(clock), .RN(n311), .Q(\U6/DATA2_4 ), 
        .QN(n247) );
  DFFR_X1 \CdfMin_reg[5]  ( .D(n449), .CK(clock), .RN(n311), .Q(\U6/DATA2_5 ), 
        .QN(n242) );
  DFFR_X1 \CdfMin_reg[6]  ( .D(n448), .CK(clock), .RN(n311), .Q(\U6/DATA2_6 ), 
        .QN(n243) );
  DFFR_X1 \CdfMin_reg[7]  ( .D(n447), .CK(clock), .RN(n311), .Q(\U6/DATA2_7 ), 
        .QN(n216) );
  DFFR_X1 \CdfMin_reg[8]  ( .D(n446), .CK(clock), .RN(n311), .Q(\U6/DATA2_8 ), 
        .QN(n228) );
  DFFR_X1 \CdfMin_reg[9]  ( .D(n445), .CK(clock), .RN(n311), .Q(\U6/DATA2_9 ), 
        .QN(n237) );
  DFFR_X1 \CdfMin_reg[10]  ( .D(n444), .CK(clock), .RN(n311), .Q(\U6/DATA2_10 ), .QN(n218) );
  DFFR_X1 \CdfMin_reg[11]  ( .D(n443), .CK(clock), .RN(n311), .Q(\U6/DATA2_11 ), .QN(n219) );
  DFFR_X1 \CdfMin_reg[12]  ( .D(n442), .CK(clock), .RN(n311), .Q(\U6/DATA2_12 ), .QN(n226) );
  DFFR_X1 \CdfMin_reg[13]  ( .D(n441), .CK(clock), .RN(n311), .Q(\U6/DATA2_13 ), .QN(n235) );
  DFFR_X1 \CdfMin_reg[14]  ( .D(n440), .CK(clock), .RN(n310), .Q(\U6/DATA2_14 ), .QN(n244) );
  DFFR_X1 \CdfMin_reg[15]  ( .D(n439), .CK(clock), .RN(n310), .Q(\U6/DATA2_15 ), .QN(n245) );
  OR3_X1 U97 ( .A1(\U6/DATA2_3 ), .A2(\U6/DATA2_4 ), .A3(\U6/DATA2_2 ), .ZN(
        n76) );
  DFFR_X2 CdfValid_reg ( .D(\U8/Z_0 ), .CK(clock), .RN(n310), .Q(CdfValid) );
  DFFR_X2 \AccumlateResult_reg[1]  ( .D(n239), .CK(clock), .RN(n310), .Q(
        \add/A[1] ), .QN(n301) );
  DFFR_X2 \AccumlateResult_reg[9]  ( .D(n231), .CK(clock), .RN(n310), .Q(
        \add/A[9] ), .QN(n272) );
  DFFR_X2 \AccumlateResult_reg[5]  ( .D(n250), .CK(clock), .RN(reset_n), .Q(
        \add/A[5] ), .QN(n298) );
  DFF_X2 \StoreAddressOut_reg[15]  ( .D(StoreAddressIn[15]), .CK(clock), .Q(
        StoreAddressOut[15]) );
  DFF_X2 \StoreAddressOut_reg[14]  ( .D(StoreAddressIn[14]), .CK(clock), .Q(
        StoreAddressOut[14]) );
  DFF_X2 \StoreAddressOut_reg[13]  ( .D(StoreAddressIn[13]), .CK(clock), .Q(
        StoreAddressOut[13]) );
  DFF_X2 \StoreAddressOut_reg[12]  ( .D(StoreAddressIn[12]), .CK(clock), .Q(
        StoreAddressOut[12]) );
  DFF_X2 \StoreAddressOut_reg[11]  ( .D(StoreAddressIn[11]), .CK(clock), .Q(
        StoreAddressOut[11]) );
  DFF_X2 \StoreAddressOut_reg[10]  ( .D(StoreAddressIn[10]), .CK(clock), .Q(
        StoreAddressOut[10]) );
  DFF_X2 \StoreAddressOut_reg[9]  ( .D(StoreAddressIn[9]), .CK(clock), .Q(
        StoreAddressOut[9]) );
  DFF_X2 \StoreAddressOut_reg[8]  ( .D(StoreAddressIn[8]), .CK(clock), .Q(
        StoreAddressOut[8]) );
  DFF_X2 \StoreAddressOut_reg[7]  ( .D(StoreAddressIn[7]), .CK(clock), .Q(
        StoreAddressOut[7]) );
  DFF_X2 \StoreAddressOut_reg[6]  ( .D(StoreAddressIn[6]), .CK(clock), .Q(
        StoreAddressOut[6]) );
  DFF_X2 \StoreAddressOut_reg[5]  ( .D(StoreAddressIn[5]), .CK(clock), .Q(
        StoreAddressOut[5]) );
  DFF_X2 \StoreAddressOut_reg[4]  ( .D(StoreAddressIn[4]), .CK(clock), .Q(
        StoreAddressOut[4]) );
  DFF_X2 \StoreAddressOut_reg[3]  ( .D(StoreAddressIn[3]), .CK(clock), .Q(
        StoreAddressOut[3]) );
  DFF_X2 \StoreAddressOut_reg[2]  ( .D(StoreAddressIn[2]), .CK(clock), .Q(
        StoreAddressOut[2]) );
  DFF_X2 \StoreAddressOut_reg[1]  ( .D(StoreAddressIn[1]), .CK(clock), .Q(
        StoreAddressOut[1]) );
  DFF_X2 \StoreAddressOut_reg[0]  ( .D(StoreAddressIn[0]), .CK(clock), .Q(
        StoreAddressOut[0]) );
  DFFR_X2 StartOut_reg ( .D(StartIn), .CK(clock), .RN(n311), .Q(StartOut) );
  DFFR_X2 \AccumlateResult_reg[19]  ( .D(n217), .CK(clock), .RN(n310), .Q(
        \add/A[19] ), .QN(n382) );
  DFFR_X2 \CdfMin_reg[19]  ( .D(n435), .CK(clock), .RN(n310), .Q(\U6/DATA2_19 ), .QN(n396) );
  DFFR_X2 \CdfMin_reg[17]  ( .D(n437), .CK(clock), .RN(n311), .Q(\U6/DATA2_17 ) );
  DFFR_X2 \CdfMin_reg[16]  ( .D(n438), .CK(clock), .RN(reset_n), .Q(
        \U6/DATA2_16 ) );
  DFFR_X2 \CdfMin_reg[18]  ( .D(n436), .CK(clock), .RN(reset_n), .Q(
        \U6/DATA2_18 ) );
  OAI221_X2 U11 ( .B1(\add/B[3] ), .B2(\add/A[3] ), .C1(n306), .C2(n260), .A(
        n325), .ZN(n332) );
  INV_X4 U15 ( .A(n358), .ZN(n258) );
  XOR2_X2 U16 ( .A(n305), .B(n389), .Z(n424) );
  NOR2_X2 U17 ( .A1(n295), .A2(n343), .ZN(n278) );
  BUF_X4 U18 ( .A(n367), .Z(n261) );
  AND4_X4 U19 ( .A1(n394), .A2(n393), .A3(n392), .A4(StartIn), .ZN(n217) );
  AND2_X4 U20 ( .A1(n288), .A2(n414), .ZN(n230) );
  AND2_X4 U21 ( .A1(StartIn), .A2(n416), .ZN(n231) );
  AND2_X4 U22 ( .A1(StartIn), .A2(n415), .ZN(n232) );
  XOR2_X2 U23 ( .A(\add/B[17] ), .B(\add/A[17] ), .Z(n233) );
  AND2_X4 U24 ( .A1(StartIn), .A2(n410), .ZN(n239) );
  AND2_X4 U25 ( .A1(StartIn), .A2(n294), .ZN(n240) );
  AND2_X1 U26 ( .A1(\U6/DATA1_5 ), .A2(StartIn), .ZN(n250) );
  INV_X2 U27 ( .A(n384), .ZN(n386) );
  NAND2_X2 U28 ( .A1(n274), .A2(n275), .ZN(n251) );
  INV_X4 U29 ( .A(n251), .ZN(n373) );
  INV_X1 U30 ( .A(n251), .ZN(n252) );
  NAND2_X1 U31 ( .A1(\add/B[1] ), .A2(n300), .ZN(n323) );
  INV_X4 U32 ( .A(n253), .ZN(n254) );
  OR3_X4 U33 ( .A1(n278), .A2(n277), .A3(n279), .ZN(n344) );
  INV_X4 U34 ( .A(n322), .ZN(n255) );
  NAND2_X1 U35 ( .A1(\add/B[3] ), .A2(\add/A[3] ), .ZN(n333) );
  NOR2_X4 U36 ( .A1(n351), .A2(n271), .ZN(n265) );
  NAND2_X2 U37 ( .A1(\add/B[2] ), .A2(\add/A[2] ), .ZN(n324) );
  AND2_X4 U38 ( .A1(n422), .A2(n421), .ZN(n305) );
  NAND2_X2 U39 ( .A1(StartIn), .A2(n425), .ZN(n256) );
  INV_X1 U40 ( .A(\add/B[2] ), .ZN(n317) );
  XNOR2_X2 U41 ( .A(n233), .B(n308), .ZN(n408) );
  NAND2_X1 U42 ( .A1(n319), .A2(n324), .ZN(n321) );
  INV_X2 U43 ( .A(n381), .ZN(n378) );
  OAI21_X4 U44 ( .B1(n381), .B2(n380), .A(n379), .ZN(n384) );
  OAI22_X1 U45 ( .A1(n281), .A2(n252), .B1(n225), .B2(n372), .ZN(n257) );
  INV_X4 U46 ( .A(n258), .ZN(n259) );
  NAND2_X2 U47 ( .A1(n324), .A2(n323), .ZN(n260) );
  NAND2_X1 U48 ( .A1(n324), .A2(n323), .ZN(n326) );
  AOI22_X2 U49 ( .A1(n347), .A2(n348), .B1(\add/B[8] ), .B2(\add/A[8] ), .ZN(
        n351) );
  AND2_X2 U50 ( .A1(n315), .A2(n301), .ZN(n307) );
  NOR2_X2 U51 ( .A1(n313), .A2(n307), .ZN(n306) );
  INV_X1 U52 ( .A(n351), .ZN(n262) );
  INV_X4 U53 ( .A(n262), .ZN(n263) );
  OAI22_X2 U54 ( .A1(n268), .A2(n367), .B1(n366), .B2(n221), .ZN(n264) );
  OAI22_X1 U55 ( .A1(n268), .A2(n261), .B1(n366), .B2(n221), .ZN(n267) );
  NOR2_X2 U56 ( .A1(n350), .A2(n272), .ZN(n266) );
  OR2_X4 U57 ( .A1(n265), .A2(n266), .ZN(n270) );
  AOI22_X2 U58 ( .A1(n270), .A2(n355), .B1(\add/B[10] ), .B2(\add/A[10] ), 
        .ZN(n358) );
  AND2_X4 U59 ( .A1(n221), .A2(n366), .ZN(n268) );
  AOI22_X2 U60 ( .A1(n364), .A2(n363), .B1(\add/B[12] ), .B2(\add/A[12] ), 
        .ZN(n367) );
  OAI22_X1 U61 ( .A1(n263), .A2(n271), .B1(n350), .B2(n272), .ZN(n269) );
  NAND2_X2 U62 ( .A1(\add/B[14] ), .A2(\add/A[14] ), .ZN(n275) );
  NAND2_X2 U63 ( .A1(n227), .A2(n369), .ZN(n370) );
  INV_X4 U64 ( .A(n269), .ZN(n354) );
  AND2_X4 U65 ( .A1(n272), .A2(n350), .ZN(n271) );
  INV_X1 U66 ( .A(n267), .ZN(n273) );
  INV_X2 U67 ( .A(\add/B[5] ), .ZN(n296) );
  NAND2_X2 U68 ( .A1(n264), .A2(n370), .ZN(n274) );
  XOR2_X1 U69 ( .A(n371), .B(n252), .Z(\U6/DATA1_15 ) );
  OAI221_X1 U70 ( .B1(\add/B[3] ), .B2(\add/A[3] ), .C1(n255), .C2(n326), .A(
        n325), .ZN(n276) );
  INV_X1 U71 ( .A(n257), .ZN(n376) );
  NOR2_X2 U72 ( .A1(\add/B[7] ), .A2(\add/A[7] ), .ZN(n277) );
  INV_X1 U73 ( .A(n342), .ZN(n279) );
  OR2_X1 U74 ( .A1(\add/A[6] ), .A2(\add/B[6] ), .ZN(n342) );
  NAND2_X1 U75 ( .A1(n387), .A2(n386), .ZN(n283) );
  AND2_X4 U76 ( .A1(n408), .A2(StartIn), .ZN(n286) );
  OR2_X2 U77 ( .A1(\add/A[8] ), .A2(\add/B[8] ), .ZN(n348) );
  XOR2_X1 U78 ( .A(n346), .B(n347), .Z(n415) );
  XNOR2_X1 U79 ( .A(\add/B[7] ), .B(\add/A[7] ), .ZN(n290) );
  XNOR2_X1 U80 ( .A(\add/B[4] ), .B(\add/A[4] ), .ZN(n291) );
  XOR2_X1 U81 ( .A(\add/A[0] ), .B(\add/B[0] ), .Z(n294) );
  XNOR2_X1 U82 ( .A(\add/B[6] ), .B(\add/A[6] ), .ZN(n292) );
  XNOR2_X1 U83 ( .A(\add/B[5] ), .B(\add/A[5] ), .ZN(n293) );
  XOR2_X1 U84 ( .A(n314), .B(n313), .Z(n410) );
  OAI22_X2 U85 ( .A1(n373), .A2(n281), .B1(n225), .B2(n372), .ZN(n280) );
  AND2_X4 U86 ( .A1(n225), .A2(n372), .ZN(n281) );
  AOI221_X1 U87 ( .B1(n296), .B2(n298), .C1(n276), .C2(n299), .A(n297), .ZN(
        n282) );
  INV_X4 U88 ( .A(n312), .ZN(n310) );
  INV_X4 U89 ( .A(n312), .ZN(n311) );
  INV_X4 U90 ( .A(reset_n), .ZN(n312) );
  AND2_X1 U91 ( .A1(n283), .A2(n284), .ZN(n394) );
  NAND2_X2 U92 ( .A1(n385), .A2(n423), .ZN(n284) );
  NAND2_X2 U93 ( .A1(StartIn), .A2(n432), .ZN(n433) );
  NOR2_X2 U94 ( .A1(n423), .A2(n391), .ZN(n387) );
  OR2_X1 U95 ( .A1(n428), .A2(n309), .ZN(n285) );
  AND2_X1 U96 ( .A1(StartIn), .A2(n409), .ZN(n287) );
  AND2_X1 U98 ( .A1(n412), .A2(n413), .ZN(n288) );
  NAND2_X2 U99 ( .A1(StartIn), .A2(n428), .ZN(n432) );
  XNOR2_X2 U100 ( .A(\add/A[13] ), .B(\add/B[13] ), .ZN(n365) );
  XNOR2_X2 U101 ( .A(\add/A[12] ), .B(\add/B[12] ), .ZN(n360) );
  XNOR2_X2 U102 ( .A(\add/A[11] ), .B(\add/B[11] ), .ZN(n356) );
  INV_X4 U103 ( .A(n335), .ZN(n297) );
  XNOR2_X2 U104 ( .A(\add/A[14] ), .B(\add/B[14] ), .ZN(n368) );
  XOR2_X2 U105 ( .A(n289), .B(n386), .Z(n425) );
  XNOR2_X2 U106 ( .A(\add/B[18] ), .B(\add/A[18] ), .ZN(n289) );
  XOR2_X2 U107 ( .A(n374), .B(n376), .Z(n409) );
  XNOR2_X2 U108 ( .A(\add/A[10] ), .B(\add/B[10] ), .ZN(n352) );
  XNOR2_X2 U109 ( .A(\add/A[9] ), .B(\add/B[9] ), .ZN(n349) );
  XNOR2_X2 U110 ( .A(n338), .B(n290), .ZN(\U6/DATA1_7 ) );
  XNOR2_X2 U111 ( .A(n329), .B(n291), .ZN(\U6/DATA1_4 ) );
  XNOR2_X2 U112 ( .A(n336), .B(n292), .ZN(\U6/DATA1_6 ) );
  XNOR2_X2 U113 ( .A(n331), .B(n293), .ZN(\U6/DATA1_5 ) );
  XOR2_X1 U114 ( .A(\add/B[3] ), .B(\add/A[3] ), .Z(n320) );
  AOI221_X2 U115 ( .B1(n298), .B2(n296), .C1(n332), .C2(n299), .A(n297), .ZN(
        n295) );
  INV_X4 U116 ( .A(n282), .ZN(n339) );
  AND2_X4 U117 ( .A1(n334), .A2(n333), .ZN(n299) );
  INV_X2 U118 ( .A(n301), .ZN(n300) );
  NAND2_X2 U119 ( .A1(n230), .A2(n411), .ZN(n427) );
  INV_X2 U120 ( .A(n256), .ZN(n302) );
  INV_X2 U121 ( .A(n421), .ZN(n385) );
  NAND2_X2 U122 ( .A1(n217), .A2(n432), .ZN(n303) );
  NAND2_X2 U123 ( .A1(\U6/DATA2_19 ), .A2(n407), .ZN(n304) );
  NAND2_X2 U124 ( .A1(n303), .A2(n304), .ZN(n435) );
  XNOR2_X1 U125 ( .A(\add/B[2] ), .B(\add/A[2] ), .ZN(n316) );
  INV_X1 U126 ( .A(n306), .ZN(n322) );
  INV_X4 U127 ( .A(n378), .ZN(n308) );
  INV_X2 U128 ( .A(\U6/DATA1_15 ), .ZN(n414) );
  INV_X1 U129 ( .A(\U6/DATA1_14 ), .ZN(n413) );
  NAND2_X1 U130 ( .A1(n323), .A2(n322), .ZN(n318) );
  NOR2_X2 U131 ( .A1(n429), .A2(n285), .ZN(\U8/Z_0 ) );
  INV_X2 U132 ( .A(\add/B[1] ), .ZN(n315) );
  INV_X4 U133 ( .A(StartIn), .ZN(n309) );
  XNOR2_X1 U134 ( .A(\add/B[1] ), .B(\add/A[1] ), .ZN(n314) );
  XOR2_X1 U135 ( .A(n365), .B(n261), .Z(\U6/DATA1_13 ) );
  XOR2_X1 U136 ( .A(n349), .B(n263), .Z(n416) );
  XOR2_X1 U137 ( .A(n368), .B(n273), .Z(\U6/DATA1_14 ) );
  XOR2_X1 U138 ( .A(n352), .B(n354), .Z(\U6/DATA1_10 ) );
  XOR2_X1 U139 ( .A(n356), .B(n259), .Z(\U6/DATA1_11 ) );
  XOR2_X1 U140 ( .A(n360), .B(n362), .Z(\U6/DATA1_12 ) );
  NAND2_X1 U141 ( .A1(n333), .A2(n276), .ZN(n329) );
  NAND2_X1 U142 ( .A1(n340), .A2(n339), .ZN(n336) );
  NAND2_X2 U143 ( .A1(\add/B[0] ), .A2(n254), .ZN(n313) );
  XNOR2_X2 U144 ( .A(n316), .B(n318), .ZN(\U6/DATA1_2 ) );
  NAND2_X2 U145 ( .A1(n220), .A2(n317), .ZN(n325) );
  NAND2_X2 U146 ( .A1(n318), .A2(n325), .ZN(n319) );
  XOR2_X2 U147 ( .A(n321), .B(n320), .Z(\U6/DATA1_3 ) );
  INV_X4 U148 ( .A(\add/A[4] ), .ZN(n328) );
  INV_X4 U149 ( .A(\add/B[4] ), .ZN(n327) );
  NAND2_X2 U150 ( .A1(n328), .A2(n327), .ZN(n335) );
  NAND2_X2 U151 ( .A1(n335), .A2(n329), .ZN(n330) );
  NAND2_X2 U152 ( .A1(\add/B[4] ), .A2(\add/A[4] ), .ZN(n334) );
  NAND2_X2 U153 ( .A1(n330), .A2(n334), .ZN(n331) );
  NAND2_X2 U154 ( .A1(\add/B[5] ), .A2(\add/A[5] ), .ZN(n340) );
  NAND2_X2 U155 ( .A1(n336), .A2(n342), .ZN(n337) );
  NAND2_X2 U156 ( .A1(\add/B[6] ), .A2(\add/A[6] ), .ZN(n341) );
  NAND2_X2 U157 ( .A1(n337), .A2(n341), .ZN(n338) );
  XOR2_X2 U158 ( .A(\add/A[8] ), .B(\add/B[8] ), .Z(n346) );
  NAND2_X2 U159 ( .A1(\add/B[7] ), .A2(\add/A[7] ), .ZN(n345) );
  NAND2_X2 U160 ( .A1(n341), .A2(n340), .ZN(n343) );
  NAND2_X2 U161 ( .A1(n345), .A2(n344), .ZN(n347) );
  INV_X4 U162 ( .A(\add/B[9] ), .ZN(n350) );
  INV_X4 U163 ( .A(\add/B[10] ), .ZN(n353) );
  NAND2_X2 U164 ( .A1(n223), .A2(n353), .ZN(n355) );
  INV_X4 U165 ( .A(\add/B[11] ), .ZN(n357) );
  NAND2_X2 U166 ( .A1(n222), .A2(n357), .ZN(n359) );
  AOI22_X4 U167 ( .A1(n258), .A2(n359), .B1(\add/B[11] ), .B2(\add/A[11] ), 
        .ZN(n362) );
  INV_X4 U168 ( .A(\add/B[12] ), .ZN(n361) );
  NAND2_X2 U169 ( .A1(n224), .A2(n361), .ZN(n364) );
  INV_X4 U170 ( .A(n362), .ZN(n363) );
  INV_X4 U171 ( .A(\add/B[13] ), .ZN(n366) );
  XNOR2_X2 U172 ( .A(\add/B[15] ), .B(\add/A[15] ), .ZN(n371) );
  INV_X4 U173 ( .A(\add/B[14] ), .ZN(n369) );
  XNOR2_X2 U174 ( .A(\add/B[16] ), .B(\add/A[16] ), .ZN(n374) );
  INV_X4 U175 ( .A(\add/B[15] ), .ZN(n372) );
  INV_X4 U176 ( .A(\add/B[16] ), .ZN(n375) );
  NAND2_X2 U177 ( .A1(n234), .A2(n375), .ZN(n377) );
  AOI22_X4 U178 ( .A1(n280), .A2(n377), .B1(\add/A[16] ), .B2(\add/B[16] ), 
        .ZN(n381) );
  NOR2_X2 U179 ( .A1(\add/B[17] ), .A2(\add/A[17] ), .ZN(n380) );
  NAND2_X2 U180 ( .A1(\add/A[17] ), .A2(\add/B[17] ), .ZN(n379) );
  XOR2_X2 U181 ( .A(n382), .B(\add/B[19] ), .Z(n389) );
  INV_X4 U182 ( .A(n389), .ZN(n423) );
  NAND2_X2 U183 ( .A1(\add/B[18] ), .A2(\add/A[18] ), .ZN(n422) );
  INV_X4 U184 ( .A(n422), .ZN(n391) );
  INV_X4 U185 ( .A(\add/B[18] ), .ZN(n383) );
  NAND2_X2 U186 ( .A1(n236), .A2(n383), .ZN(n388) );
  NAND2_X2 U187 ( .A1(n384), .A2(n388), .ZN(n421) );
  INV_X4 U188 ( .A(n388), .ZN(n390) );
  NAND2_X2 U189 ( .A1(n390), .A2(n389), .ZN(n393) );
  NAND2_X2 U190 ( .A1(n391), .A2(n423), .ZN(n392) );
  NAND3_X2 U191 ( .A1(n219), .A2(n226), .A3(n235), .ZN(n395) );
  NOR3_X2 U192 ( .A1(n395), .A2(\U6/DATA2_15 ), .A3(\U6/DATA2_14 ), .ZN(n401)
         );
  NOR4_X2 U193 ( .A1(n76), .A2(\U6/DATA2_18 ), .A3(\U6/DATA2_17 ), .A4(
        \U6/DATA2_16 ), .ZN(n400) );
  NAND4_X2 U194 ( .A1(n216), .A2(n228), .A3(n237), .A4(n218), .ZN(n398) );
  NAND3_X2 U195 ( .A1(n396), .A2(n229), .A3(n238), .ZN(n397) );
  NOR4_X2 U196 ( .A1(n398), .A2(n397), .A3(\U6/DATA2_6 ), .A4(\U6/DATA2_5 ), 
        .ZN(n399) );
  NAND3_X2 U197 ( .A1(n401), .A2(n400), .A3(n399), .ZN(n428) );
  INV_X4 U198 ( .A(n432), .ZN(n407) );
  MUX2_X2 U199 ( .A(n240), .B(\U6/DATA2_0 ), .S(n407), .Z(n454) );
  MUX2_X2 U200 ( .A(n239), .B(\U6/DATA2_1 ), .S(n407), .Z(n453) );
  INV_X4 U201 ( .A(\U6/DATA1_5 ), .ZN(n419) );
  OAI22_X2 U202 ( .A1(n419), .A2(n433), .B1(n432), .B2(n242), .ZN(n449) );
  INV_X4 U203 ( .A(\U6/DATA1_6 ), .ZN(n420) );
  OAI22_X2 U204 ( .A1(n420), .A2(n433), .B1(n432), .B2(n243), .ZN(n448) );
  INV_X4 U205 ( .A(\U6/DATA1_7 ), .ZN(n402) );
  OAI22_X2 U206 ( .A1(n402), .A2(n433), .B1(n432), .B2(n216), .ZN(n447) );
  MUX2_X2 U207 ( .A(n232), .B(\U6/DATA2_8 ), .S(n407), .Z(n446) );
  MUX2_X2 U208 ( .A(n231), .B(\U6/DATA2_9 ), .S(n407), .Z(n445) );
  INV_X4 U209 ( .A(\U6/DATA1_10 ), .ZN(n403) );
  OAI22_X2 U210 ( .A1(n403), .A2(n433), .B1(n432), .B2(n218), .ZN(n444) );
  INV_X4 U211 ( .A(\U6/DATA1_11 ), .ZN(n404) );
  OAI22_X2 U212 ( .A1(n404), .A2(n433), .B1(n432), .B2(n219), .ZN(n443) );
  INV_X4 U213 ( .A(\U6/DATA1_12 ), .ZN(n405) );
  OAI22_X2 U214 ( .A1(n405), .A2(n433), .B1(n432), .B2(n226), .ZN(n442) );
  INV_X4 U215 ( .A(\U6/DATA1_13 ), .ZN(n406) );
  OAI22_X2 U216 ( .A1(n406), .A2(n433), .B1(n432), .B2(n235), .ZN(n441) );
  OAI22_X2 U217 ( .A1(n413), .A2(n433), .B1(n432), .B2(n244), .ZN(n440) );
  OAI22_X2 U218 ( .A1(n414), .A2(n433), .B1(n432), .B2(n245), .ZN(n439) );
  MUX2_X2 U219 ( .A(n287), .B(\U6/DATA2_16 ), .S(n407), .Z(n438) );
  MUX2_X2 U220 ( .A(n286), .B(\U6/DATA2_17 ), .S(n407), .Z(n437) );
  MUX2_X2 U221 ( .A(n302), .B(\U6/DATA2_18 ), .S(n407), .Z(n436) );
  NOR3_X2 U222 ( .A1(\U6/DATA1_13 ), .A2(\U6/DATA1_11 ), .A3(\U6/DATA1_12 ), 
        .ZN(n412) );
  NOR4_X2 U223 ( .A1(n410), .A2(n408), .A3(n409), .A4(n294), .ZN(n411) );
  NOR3_X2 U224 ( .A1(\U6/DATA1_4 ), .A2(\U6/DATA1_3 ), .A3(\U6/DATA1_2 ), .ZN(
        n418) );
  NOR4_X2 U225 ( .A1(n416), .A2(\U6/DATA1_10 ), .A3(\U6/DATA1_7 ), .A4(n415), 
        .ZN(n417) );
  NAND4_X2 U226 ( .A1(n420), .A2(n419), .A3(n418), .A4(n417), .ZN(n426) );
  NOR4_X2 U227 ( .A1(n427), .A2(n426), .A3(n425), .A4(n424), .ZN(n429) );
  INV_X4 U228 ( .A(\U6/DATA1_2 ), .ZN(n430) );
  OAI22_X2 U229 ( .A1(n430), .A2(n433), .B1(n432), .B2(n248), .ZN(n452) );
  INV_X4 U230 ( .A(\U6/DATA1_3 ), .ZN(n431) );
  OAI22_X2 U231 ( .A1(n431), .A2(n433), .B1(n432), .B2(n246), .ZN(n451) );
  INV_X4 U232 ( .A(\U6/DATA1_4 ), .ZN(n434) );
  OAI22_X2 U233 ( .A1(n434), .A2(n433), .B1(n432), .B2(n247), .ZN(n450) );
endmodule


module Cdf_Store ( clock, reset_n, StartIn, ResultIn, StoreAddressIn, WriteBus, 
        WriteAddress, WriteEnable );
  input [19:0] ResultIn;
  input [15:0] StoreAddressIn;
  output [127:0] WriteBus;
  output [15:0] WriteAddress;
  input clock, reset_n, StartIn;
  output WriteEnable;
  wire   \U5/Z_0 , \U5/Z_1 , \U5/Z_2 , \U5/Z_3 , \U5/Z_4 , \U5/Z_5 , \U5/Z_6 ,
         \U5/Z_7 , \U5/Z_8 , \U5/Z_9 , \U5/Z_10 , \U5/Z_11 , \U5/Z_12 ,
         \U5/Z_13 , \U5/Z_14 , \U5/Z_15 , \U5/Z_16 , \U5/Z_17 , \U5/Z_18 ,
         \U5/Z_19 , \U5/DATA1_0 , \U5/DATA1_1 , \U5/DATA1_2 , \U5/DATA1_3 ,
         \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 , \U5/DATA1_7 , \U5/DATA1_8 ,
         \U5/DATA1_9 , \U5/DATA1_10 , \U5/DATA1_11 , \U5/DATA1_12 ,
         \U5/DATA1_13 , \U5/DATA1_14 , \U5/DATA1_15 , \U5/DATA1_16 ,
         \U5/DATA1_17 , \U5/DATA1_18 , \U5/DATA1_19 , \U4/Z_0 , \U4/Z_1 ,
         \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 , \U4/Z_7 , \U4/Z_8 ,
         \U4/Z_9 , \U4/Z_10 , \U4/Z_11 , \U4/Z_12 , \U4/Z_13 , \U4/Z_14 ,
         \U4/Z_15 , \U4/DATA1_0 , \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 ,
         \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 , \U4/DATA1_7 , \U4/DATA1_8 ,
         \U4/DATA1_9 , \U4/DATA1_10 , \U4/DATA1_11 , \U4/DATA1_12 ,
         \U4/DATA1_13 , \U4/DATA1_14 , \U4/DATA1_15 , n443, n444, n445, n446;
  assign \U5/DATA1_0  = ResultIn[0];
  assign \U5/DATA1_1  = ResultIn[1];
  assign \U5/DATA1_2  = ResultIn[2];
  assign \U5/DATA1_3  = ResultIn[3];
  assign \U5/DATA1_4  = ResultIn[4];
  assign \U5/DATA1_5  = ResultIn[5];
  assign \U5/DATA1_6  = ResultIn[6];
  assign \U5/DATA1_7  = ResultIn[7];
  assign \U5/DATA1_8  = ResultIn[8];
  assign \U5/DATA1_9  = ResultIn[9];
  assign \U5/DATA1_10  = ResultIn[10];
  assign \U5/DATA1_11  = ResultIn[11];
  assign \U5/DATA1_12  = ResultIn[12];
  assign \U5/DATA1_13  = ResultIn[13];
  assign \U5/DATA1_14  = ResultIn[14];
  assign \U5/DATA1_15  = ResultIn[15];
  assign \U5/DATA1_16  = ResultIn[16];
  assign \U5/DATA1_17  = ResultIn[17];
  assign \U5/DATA1_18  = ResultIn[18];
  assign \U5/DATA1_19  = ResultIn[19];
  assign \U4/DATA1_0  = StoreAddressIn[0];
  assign \U4/DATA1_1  = StoreAddressIn[1];
  assign \U4/DATA1_2  = StoreAddressIn[2];
  assign \U4/DATA1_3  = StoreAddressIn[3];
  assign \U4/DATA1_4  = StoreAddressIn[4];
  assign \U4/DATA1_5  = StoreAddressIn[5];
  assign \U4/DATA1_6  = StoreAddressIn[6];
  assign \U4/DATA1_7  = StoreAddressIn[7];
  assign \U4/DATA1_8  = StoreAddressIn[8];
  assign \U4/DATA1_9  = StoreAddressIn[9];
  assign \U4/DATA1_10  = StoreAddressIn[10];
  assign \U4/DATA1_11  = StoreAddressIn[11];
  assign \U4/DATA1_12  = StoreAddressIn[12];
  assign \U4/DATA1_13  = StoreAddressIn[13];
  assign \U4/DATA1_14  = StoreAddressIn[14];
  assign \U4/DATA1_15  = StoreAddressIn[15];

  DFFR_X1 \WriteBus_reg[14]  ( .D(\U5/Z_14 ), .CK(clock), .RN(n446), .Q(
        WriteBus[14]) );
  DFFR_X1 \WriteBus_reg[13]  ( .D(\U5/Z_13 ), .CK(clock), .RN(n446), .Q(
        WriteBus[13]) );
  DFFR_X1 \WriteBus_reg[12]  ( .D(\U5/Z_12 ), .CK(clock), .RN(n446), .Q(
        WriteBus[12]) );
  DFFR_X1 \WriteBus_reg[11]  ( .D(\U5/Z_11 ), .CK(clock), .RN(n446), .Q(
        WriteBus[11]) );
  DFFR_X1 \WriteBus_reg[10]  ( .D(\U5/Z_10 ), .CK(clock), .RN(n446), .Q(
        WriteBus[10]) );
  DFFR_X1 \WriteBus_reg[9]  ( .D(\U5/Z_9 ), .CK(clock), .RN(n446), .Q(
        WriteBus[9]) );
  DFFR_X1 \WriteBus_reg[8]  ( .D(\U5/Z_8 ), .CK(clock), .RN(n446), .Q(
        WriteBus[8]) );
  DFFR_X1 \WriteBus_reg[7]  ( .D(\U5/Z_7 ), .CK(clock), .RN(n446), .Q(
        WriteBus[7]) );
  DFFR_X1 \WriteBus_reg[6]  ( .D(\U5/Z_6 ), .CK(clock), .RN(n445), .Q(
        WriteBus[6]) );
  DFFR_X1 \WriteBus_reg[5]  ( .D(\U5/Z_5 ), .CK(clock), .RN(n445), .Q(
        WriteBus[5]) );
  DFFR_X1 \WriteBus_reg[4]  ( .D(\U5/Z_4 ), .CK(clock), .RN(n445), .Q(
        WriteBus[4]) );
  DFFR_X1 \WriteBus_reg[3]  ( .D(\U5/Z_3 ), .CK(clock), .RN(n445), .Q(
        WriteBus[3]) );
  DFFR_X1 \WriteBus_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .RN(n445), .Q(
        WriteBus[2]) );
  DFFR_X1 \WriteBus_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .RN(n445), .Q(
        WriteBus[1]) );
  DFFR_X1 \WriteBus_reg[0]  ( .D(\U5/Z_0 ), .CK(clock), .RN(n445), .Q(
        WriteBus[0]) );
  DFFR_X1 \WriteAddress_reg[15]  ( .D(\U4/Z_15 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[15]) );
  DFFR_X1 \WriteAddress_reg[14]  ( .D(\U4/Z_14 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[14]) );
  DFFR_X1 \WriteAddress_reg[13]  ( .D(\U4/Z_13 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[13]) );
  DFFR_X1 \WriteAddress_reg[12]  ( .D(\U4/Z_12 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[12]) );
  DFFR_X1 \WriteAddress_reg[11]  ( .D(\U4/Z_11 ), .CK(clock), .RN(n445), .Q(
        WriteAddress[11]) );
  DFFR_X1 \WriteAddress_reg[10]  ( .D(\U4/Z_10 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[10]) );
  DFFR_X1 \WriteAddress_reg[9]  ( .D(\U4/Z_9 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[9]) );
  DFFR_X1 \WriteAddress_reg[8]  ( .D(\U4/Z_8 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[8]) );
  DFFR_X1 \WriteAddress_reg[7]  ( .D(\U4/Z_7 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[7]) );
  DFFR_X1 \WriteAddress_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[6]) );
  DFFR_X1 \WriteAddress_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[5]) );
  DFFR_X1 \WriteAddress_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[4]) );
  DFFR_X1 \WriteAddress_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[3]) );
  DFFR_X1 \WriteAddress_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[2]) );
  DFFR_X1 \WriteAddress_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[1]) );
  DFFR_X1 \WriteAddress_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n444), .Q(
        WriteAddress[0]) );
  AND2_X1 U111 ( .A1(\U5/DATA1_9 ), .A2(StartIn), .ZN(\U5/Z_9 ) );
  AND2_X1 U112 ( .A1(\U5/DATA1_8 ), .A2(StartIn), .ZN(\U5/Z_8 ) );
  AND2_X1 U113 ( .A1(\U5/DATA1_7 ), .A2(StartIn), .ZN(\U5/Z_7 ) );
  AND2_X1 U114 ( .A1(\U5/DATA1_6 ), .A2(StartIn), .ZN(\U5/Z_6 ) );
  AND2_X1 U115 ( .A1(\U5/DATA1_5 ), .A2(StartIn), .ZN(\U5/Z_5 ) );
  AND2_X1 U116 ( .A1(\U5/DATA1_4 ), .A2(StartIn), .ZN(\U5/Z_4 ) );
  AND2_X1 U117 ( .A1(\U5/DATA1_3 ), .A2(StartIn), .ZN(\U5/Z_3 ) );
  AND2_X1 U118 ( .A1(\U5/DATA1_2 ), .A2(StartIn), .ZN(\U5/Z_2 ) );
  AND2_X1 U119 ( .A1(\U5/DATA1_19 ), .A2(StartIn), .ZN(\U5/Z_19 ) );
  AND2_X1 U120 ( .A1(\U5/DATA1_18 ), .A2(StartIn), .ZN(\U5/Z_18 ) );
  AND2_X1 U121 ( .A1(\U5/DATA1_17 ), .A2(StartIn), .ZN(\U5/Z_17 ) );
  AND2_X1 U122 ( .A1(\U5/DATA1_16 ), .A2(StartIn), .ZN(\U5/Z_16 ) );
  AND2_X1 U123 ( .A1(\U5/DATA1_15 ), .A2(StartIn), .ZN(\U5/Z_15 ) );
  AND2_X1 U124 ( .A1(\U5/DATA1_14 ), .A2(StartIn), .ZN(\U5/Z_14 ) );
  AND2_X1 U125 ( .A1(\U5/DATA1_13 ), .A2(StartIn), .ZN(\U5/Z_13 ) );
  AND2_X1 U126 ( .A1(\U5/DATA1_12 ), .A2(StartIn), .ZN(\U5/Z_12 ) );
  AND2_X1 U127 ( .A1(\U5/DATA1_11 ), .A2(StartIn), .ZN(\U5/Z_11 ) );
  AND2_X1 U128 ( .A1(\U5/DATA1_10 ), .A2(StartIn), .ZN(\U5/Z_10 ) );
  AND2_X1 U131 ( .A1(\U4/DATA1_9 ), .A2(StartIn), .ZN(\U4/Z_9 ) );
  AND2_X1 U132 ( .A1(\U4/DATA1_8 ), .A2(StartIn), .ZN(\U4/Z_8 ) );
  AND2_X1 U133 ( .A1(\U4/DATA1_7 ), .A2(StartIn), .ZN(\U4/Z_7 ) );
  AND2_X1 U134 ( .A1(\U4/DATA1_6 ), .A2(StartIn), .ZN(\U4/Z_6 ) );
  AND2_X1 U135 ( .A1(\U4/DATA1_5 ), .A2(StartIn), .ZN(\U4/Z_5 ) );
  AND2_X1 U136 ( .A1(\U4/DATA1_4 ), .A2(StartIn), .ZN(\U4/Z_4 ) );
  AND2_X1 U137 ( .A1(\U4/DATA1_3 ), .A2(StartIn), .ZN(\U4/Z_3 ) );
  AND2_X1 U138 ( .A1(\U4/DATA1_2 ), .A2(StartIn), .ZN(\U4/Z_2 ) );
  AND2_X1 U139 ( .A1(\U4/DATA1_15 ), .A2(StartIn), .ZN(\U4/Z_15 ) );
  AND2_X1 U140 ( .A1(\U4/DATA1_14 ), .A2(StartIn), .ZN(\U4/Z_14 ) );
  AND2_X1 U141 ( .A1(\U4/DATA1_13 ), .A2(StartIn), .ZN(\U4/Z_13 ) );
  AND2_X1 U142 ( .A1(\U4/DATA1_12 ), .A2(StartIn), .ZN(\U4/Z_12 ) );
  AND2_X1 U143 ( .A1(\U4/DATA1_11 ), .A2(StartIn), .ZN(\U4/Z_11 ) );
  AND2_X1 U144 ( .A1(\U4/DATA1_10 ), .A2(StartIn), .ZN(\U4/Z_10 ) );
  AND2_X1 U145 ( .A1(\U4/DATA1_1 ), .A2(StartIn), .ZN(\U4/Z_1 ) );
  AND2_X1 U146 ( .A1(\U4/DATA1_0 ), .A2(StartIn), .ZN(\U4/Z_0 ) );
  DFFR_X2 WriteEnable_reg ( .D(StartIn), .CK(clock), .RN(n444), .Q(WriteEnable) );
  DFFR_X2 \WriteBus_reg[19]  ( .D(\U5/Z_19 ), .CK(clock), .RN(reset_n), .Q(
        WriteBus[19]) );
  DFFR_X2 \WriteBus_reg[18]  ( .D(\U5/Z_18 ), .CK(clock), .RN(n446), .Q(
        WriteBus[18]) );
  DFFR_X2 \WriteBus_reg[17]  ( .D(\U5/Z_17 ), .CK(clock), .RN(n446), .Q(
        WriteBus[17]) );
  DFFR_X2 \WriteBus_reg[16]  ( .D(\U5/Z_16 ), .CK(clock), .RN(n446), .Q(
        WriteBus[16]) );
  DFFR_X2 \WriteBus_reg[15]  ( .D(\U5/Z_15 ), .CK(clock), .RN(n446), .Q(
        WriteBus[15]) );
  INV_X4 U129 ( .A(1'b1), .ZN(WriteBus[20]) );
  INV_X4 U147 ( .A(1'b1), .ZN(WriteBus[21]) );
  INV_X4 U149 ( .A(1'b1), .ZN(WriteBus[22]) );
  INV_X4 U151 ( .A(1'b1), .ZN(WriteBus[23]) );
  INV_X4 U153 ( .A(1'b1), .ZN(WriteBus[24]) );
  INV_X4 U155 ( .A(1'b1), .ZN(WriteBus[25]) );
  INV_X4 U157 ( .A(1'b1), .ZN(WriteBus[26]) );
  INV_X4 U159 ( .A(1'b1), .ZN(WriteBus[27]) );
  INV_X4 U161 ( .A(1'b1), .ZN(WriteBus[28]) );
  INV_X4 U163 ( .A(1'b1), .ZN(WriteBus[29]) );
  INV_X4 U165 ( .A(1'b1), .ZN(WriteBus[30]) );
  INV_X4 U167 ( .A(1'b1), .ZN(WriteBus[31]) );
  INV_X4 U169 ( .A(1'b1), .ZN(WriteBus[32]) );
  INV_X4 U171 ( .A(1'b1), .ZN(WriteBus[33]) );
  INV_X4 U173 ( .A(1'b1), .ZN(WriteBus[34]) );
  INV_X4 U175 ( .A(1'b1), .ZN(WriteBus[35]) );
  INV_X4 U177 ( .A(1'b1), .ZN(WriteBus[36]) );
  INV_X4 U179 ( .A(1'b1), .ZN(WriteBus[37]) );
  INV_X4 U181 ( .A(1'b1), .ZN(WriteBus[38]) );
  INV_X4 U183 ( .A(1'b1), .ZN(WriteBus[39]) );
  INV_X4 U185 ( .A(1'b1), .ZN(WriteBus[40]) );
  INV_X4 U187 ( .A(1'b1), .ZN(WriteBus[41]) );
  INV_X4 U189 ( .A(1'b1), .ZN(WriteBus[42]) );
  INV_X4 U191 ( .A(1'b1), .ZN(WriteBus[43]) );
  INV_X4 U193 ( .A(1'b1), .ZN(WriteBus[44]) );
  INV_X4 U195 ( .A(1'b1), .ZN(WriteBus[45]) );
  INV_X4 U197 ( .A(1'b1), .ZN(WriteBus[46]) );
  INV_X4 U199 ( .A(1'b1), .ZN(WriteBus[47]) );
  INV_X4 U201 ( .A(1'b1), .ZN(WriteBus[48]) );
  INV_X4 U203 ( .A(1'b1), .ZN(WriteBus[49]) );
  INV_X4 U205 ( .A(1'b1), .ZN(WriteBus[50]) );
  INV_X4 U207 ( .A(1'b1), .ZN(WriteBus[51]) );
  INV_X4 U209 ( .A(1'b1), .ZN(WriteBus[52]) );
  INV_X4 U211 ( .A(1'b1), .ZN(WriteBus[53]) );
  INV_X4 U213 ( .A(1'b1), .ZN(WriteBus[54]) );
  INV_X4 U215 ( .A(1'b1), .ZN(WriteBus[55]) );
  INV_X4 U217 ( .A(1'b1), .ZN(WriteBus[56]) );
  INV_X4 U219 ( .A(1'b1), .ZN(WriteBus[57]) );
  INV_X4 U221 ( .A(1'b1), .ZN(WriteBus[58]) );
  INV_X4 U223 ( .A(1'b1), .ZN(WriteBus[59]) );
  INV_X4 U225 ( .A(1'b1), .ZN(WriteBus[60]) );
  INV_X4 U227 ( .A(1'b1), .ZN(WriteBus[61]) );
  INV_X4 U229 ( .A(1'b1), .ZN(WriteBus[62]) );
  INV_X4 U231 ( .A(1'b1), .ZN(WriteBus[63]) );
  INV_X4 U233 ( .A(1'b1), .ZN(WriteBus[64]) );
  INV_X4 U235 ( .A(1'b1), .ZN(WriteBus[65]) );
  INV_X4 U237 ( .A(1'b1), .ZN(WriteBus[66]) );
  INV_X4 U239 ( .A(1'b1), .ZN(WriteBus[67]) );
  INV_X4 U241 ( .A(1'b1), .ZN(WriteBus[68]) );
  INV_X4 U243 ( .A(1'b1), .ZN(WriteBus[69]) );
  INV_X4 U245 ( .A(1'b1), .ZN(WriteBus[70]) );
  INV_X4 U247 ( .A(1'b1), .ZN(WriteBus[71]) );
  INV_X4 U249 ( .A(1'b1), .ZN(WriteBus[72]) );
  INV_X4 U251 ( .A(1'b1), .ZN(WriteBus[73]) );
  INV_X4 U253 ( .A(1'b1), .ZN(WriteBus[74]) );
  INV_X4 U255 ( .A(1'b1), .ZN(WriteBus[75]) );
  INV_X4 U257 ( .A(1'b1), .ZN(WriteBus[76]) );
  INV_X4 U259 ( .A(1'b1), .ZN(WriteBus[77]) );
  INV_X4 U261 ( .A(1'b1), .ZN(WriteBus[78]) );
  INV_X4 U263 ( .A(1'b1), .ZN(WriteBus[79]) );
  INV_X4 U265 ( .A(1'b1), .ZN(WriteBus[80]) );
  INV_X4 U267 ( .A(1'b1), .ZN(WriteBus[81]) );
  INV_X4 U269 ( .A(1'b1), .ZN(WriteBus[82]) );
  INV_X4 U271 ( .A(1'b1), .ZN(WriteBus[83]) );
  INV_X4 U273 ( .A(1'b1), .ZN(WriteBus[84]) );
  INV_X4 U275 ( .A(1'b1), .ZN(WriteBus[85]) );
  INV_X4 U277 ( .A(1'b1), .ZN(WriteBus[86]) );
  INV_X4 U279 ( .A(1'b1), .ZN(WriteBus[87]) );
  INV_X4 U281 ( .A(1'b1), .ZN(WriteBus[88]) );
  INV_X4 U283 ( .A(1'b1), .ZN(WriteBus[89]) );
  INV_X4 U285 ( .A(1'b1), .ZN(WriteBus[90]) );
  INV_X4 U287 ( .A(1'b1), .ZN(WriteBus[91]) );
  INV_X4 U289 ( .A(1'b1), .ZN(WriteBus[92]) );
  INV_X4 U291 ( .A(1'b1), .ZN(WriteBus[93]) );
  INV_X4 U293 ( .A(1'b1), .ZN(WriteBus[94]) );
  INV_X4 U295 ( .A(1'b1), .ZN(WriteBus[95]) );
  INV_X4 U297 ( .A(1'b1), .ZN(WriteBus[96]) );
  INV_X4 U299 ( .A(1'b1), .ZN(WriteBus[97]) );
  INV_X4 U301 ( .A(1'b1), .ZN(WriteBus[98]) );
  INV_X4 U303 ( .A(1'b1), .ZN(WriteBus[99]) );
  INV_X4 U305 ( .A(1'b1), .ZN(WriteBus[100]) );
  INV_X4 U307 ( .A(1'b1), .ZN(WriteBus[101]) );
  INV_X4 U309 ( .A(1'b1), .ZN(WriteBus[102]) );
  INV_X4 U311 ( .A(1'b1), .ZN(WriteBus[103]) );
  INV_X4 U313 ( .A(1'b1), .ZN(WriteBus[104]) );
  INV_X4 U315 ( .A(1'b1), .ZN(WriteBus[105]) );
  INV_X4 U317 ( .A(1'b1), .ZN(WriteBus[106]) );
  INV_X4 U319 ( .A(1'b1), .ZN(WriteBus[107]) );
  INV_X4 U321 ( .A(1'b1), .ZN(WriteBus[108]) );
  INV_X4 U323 ( .A(1'b1), .ZN(WriteBus[109]) );
  INV_X4 U325 ( .A(1'b1), .ZN(WriteBus[110]) );
  INV_X4 U327 ( .A(1'b1), .ZN(WriteBus[111]) );
  INV_X4 U329 ( .A(1'b1), .ZN(WriteBus[112]) );
  INV_X4 U331 ( .A(1'b1), .ZN(WriteBus[113]) );
  INV_X4 U333 ( .A(1'b1), .ZN(WriteBus[114]) );
  INV_X4 U335 ( .A(1'b1), .ZN(WriteBus[115]) );
  INV_X4 U337 ( .A(1'b1), .ZN(WriteBus[116]) );
  INV_X4 U339 ( .A(1'b1), .ZN(WriteBus[117]) );
  INV_X4 U341 ( .A(1'b1), .ZN(WriteBus[118]) );
  INV_X4 U343 ( .A(1'b1), .ZN(WriteBus[119]) );
  INV_X4 U345 ( .A(1'b1), .ZN(WriteBus[120]) );
  INV_X4 U347 ( .A(1'b1), .ZN(WriteBus[121]) );
  INV_X4 U349 ( .A(1'b1), .ZN(WriteBus[122]) );
  INV_X4 U351 ( .A(1'b1), .ZN(WriteBus[123]) );
  INV_X4 U353 ( .A(1'b1), .ZN(WriteBus[124]) );
  INV_X4 U355 ( .A(1'b1), .ZN(WriteBus[125]) );
  INV_X4 U357 ( .A(1'b1), .ZN(WriteBus[126]) );
  INV_X4 U359 ( .A(1'b1), .ZN(WriteBus[127]) );
  INV_X4 U361 ( .A(n443), .ZN(n445) );
  INV_X4 U362 ( .A(n443), .ZN(n446) );
  INV_X4 U363 ( .A(n443), .ZN(n444) );
  INV_X4 U364 ( .A(reset_n), .ZN(n443) );
  AND2_X4 U365 ( .A1(\U5/DATA1_1 ), .A2(StartIn), .ZN(\U5/Z_1 ) );
  AND2_X4 U366 ( .A1(\U5/DATA1_0 ), .A2(StartIn), .ZN(\U5/Z_0 ) );
endmodule


module Cdf_top ( clock, reset_n, start, SP_ReadBus, SP_ReadAddress, 
        WriteEnable, Output_MEMBus, Output_MEMAddress, Cdf_Min, done, 
        input_base_offset, cdf_valid );
  input [35:0] SP_ReadBus;
  output [15:0] SP_ReadAddress;
  output [127:0] Output_MEMBus;
  output [15:0] Output_MEMAddress;
  output [19:0] Cdf_Min;
  input clock, reset_n, start, input_base_offset;
  output WriteEnable, done, cdf_valid;
  wire   start_to_accumlate, start_to_store, n217, n218;
  wire   [19:0] Accumlate;
  wire   [19:0] AccumlateResult;
  wire   [15:0] store_address;
  wire   [15:0] store_address_to_store;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107;

  Cdf_Fetch stage1 ( .clock(clock), .reset_n(n217), .start(start), .ReadBus(
        SP_ReadBus), .ReadAddr(SP_ReadAddress), .AccumlateOut(Accumlate), 
        .StartOut(start_to_accumlate), .StoreAddress(store_address), 
        .input_base_offset(input_base_offset), .done(done) );
  Cdf_Accumlate stage2 ( .clock(clock), .reset_n(n217), .AccumlateIn(Accumlate), .StartIn(start_to_accumlate), .StoreAddressIn(store_address), 
        .AccumlateResult(AccumlateResult), .StoreAddressOut(
        store_address_to_store), .StartOut(start_to_store), .CdfMin(Cdf_Min), 
        .CdfValid(cdf_valid) );
  Cdf_Store stage3 ( .clock(clock), .reset_n(n217), .StartIn(start_to_store), 
        .ResultIn(AccumlateResult), .StoreAddressIn(store_address_to_store), 
        .WriteBus({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        Output_MEMBus[19:0]}), .WriteAddress(Output_MEMAddress), .WriteEnable(
        WriteEnable) );
  INV_X4 U1 ( .A(1'b1), .ZN(Output_MEMBus[20]) );
  INV_X4 U3 ( .A(1'b1), .ZN(Output_MEMBus[21]) );
  INV_X4 U5 ( .A(1'b1), .ZN(Output_MEMBus[22]) );
  INV_X4 U7 ( .A(1'b1), .ZN(Output_MEMBus[23]) );
  INV_X4 U9 ( .A(1'b1), .ZN(Output_MEMBus[24]) );
  INV_X4 U11 ( .A(1'b1), .ZN(Output_MEMBus[25]) );
  INV_X4 U13 ( .A(1'b1), .ZN(Output_MEMBus[26]) );
  INV_X4 U15 ( .A(1'b1), .ZN(Output_MEMBus[27]) );
  INV_X4 U17 ( .A(1'b1), .ZN(Output_MEMBus[28]) );
  INV_X4 U19 ( .A(1'b1), .ZN(Output_MEMBus[29]) );
  INV_X4 U21 ( .A(1'b1), .ZN(Output_MEMBus[30]) );
  INV_X4 U23 ( .A(1'b1), .ZN(Output_MEMBus[31]) );
  INV_X4 U25 ( .A(1'b1), .ZN(Output_MEMBus[32]) );
  INV_X4 U27 ( .A(1'b1), .ZN(Output_MEMBus[33]) );
  INV_X4 U29 ( .A(1'b1), .ZN(Output_MEMBus[34]) );
  INV_X4 U31 ( .A(1'b1), .ZN(Output_MEMBus[35]) );
  INV_X4 U33 ( .A(1'b1), .ZN(Output_MEMBus[36]) );
  INV_X4 U35 ( .A(1'b1), .ZN(Output_MEMBus[37]) );
  INV_X4 U37 ( .A(1'b1), .ZN(Output_MEMBus[38]) );
  INV_X4 U39 ( .A(1'b1), .ZN(Output_MEMBus[39]) );
  INV_X4 U41 ( .A(1'b1), .ZN(Output_MEMBus[40]) );
  INV_X4 U43 ( .A(1'b1), .ZN(Output_MEMBus[41]) );
  INV_X4 U45 ( .A(1'b1), .ZN(Output_MEMBus[42]) );
  INV_X4 U47 ( .A(1'b1), .ZN(Output_MEMBus[43]) );
  INV_X4 U49 ( .A(1'b1), .ZN(Output_MEMBus[44]) );
  INV_X4 U51 ( .A(1'b1), .ZN(Output_MEMBus[45]) );
  INV_X4 U53 ( .A(1'b1), .ZN(Output_MEMBus[46]) );
  INV_X4 U55 ( .A(1'b1), .ZN(Output_MEMBus[47]) );
  INV_X4 U57 ( .A(1'b1), .ZN(Output_MEMBus[48]) );
  INV_X4 U59 ( .A(1'b1), .ZN(Output_MEMBus[49]) );
  INV_X4 U61 ( .A(1'b1), .ZN(Output_MEMBus[50]) );
  INV_X4 U63 ( .A(1'b1), .ZN(Output_MEMBus[51]) );
  INV_X4 U65 ( .A(1'b1), .ZN(Output_MEMBus[52]) );
  INV_X4 U67 ( .A(1'b1), .ZN(Output_MEMBus[53]) );
  INV_X4 U69 ( .A(1'b1), .ZN(Output_MEMBus[54]) );
  INV_X4 U71 ( .A(1'b1), .ZN(Output_MEMBus[55]) );
  INV_X4 U73 ( .A(1'b1), .ZN(Output_MEMBus[56]) );
  INV_X4 U75 ( .A(1'b1), .ZN(Output_MEMBus[57]) );
  INV_X4 U77 ( .A(1'b1), .ZN(Output_MEMBus[58]) );
  INV_X4 U79 ( .A(1'b1), .ZN(Output_MEMBus[59]) );
  INV_X4 U81 ( .A(1'b1), .ZN(Output_MEMBus[60]) );
  INV_X4 U83 ( .A(1'b1), .ZN(Output_MEMBus[61]) );
  INV_X4 U85 ( .A(1'b1), .ZN(Output_MEMBus[62]) );
  INV_X4 U87 ( .A(1'b1), .ZN(Output_MEMBus[63]) );
  INV_X4 U89 ( .A(1'b1), .ZN(Output_MEMBus[64]) );
  INV_X4 U91 ( .A(1'b1), .ZN(Output_MEMBus[65]) );
  INV_X4 U93 ( .A(1'b1), .ZN(Output_MEMBus[66]) );
  INV_X4 U95 ( .A(1'b1), .ZN(Output_MEMBus[67]) );
  INV_X4 U97 ( .A(1'b1), .ZN(Output_MEMBus[68]) );
  INV_X4 U99 ( .A(1'b1), .ZN(Output_MEMBus[69]) );
  INV_X4 U101 ( .A(1'b1), .ZN(Output_MEMBus[70]) );
  INV_X4 U103 ( .A(1'b1), .ZN(Output_MEMBus[71]) );
  INV_X4 U105 ( .A(1'b1), .ZN(Output_MEMBus[72]) );
  INV_X4 U107 ( .A(1'b1), .ZN(Output_MEMBus[73]) );
  INV_X4 U109 ( .A(1'b1), .ZN(Output_MEMBus[74]) );
  INV_X4 U111 ( .A(1'b1), .ZN(Output_MEMBus[75]) );
  INV_X4 U113 ( .A(1'b1), .ZN(Output_MEMBus[76]) );
  INV_X4 U115 ( .A(1'b1), .ZN(Output_MEMBus[77]) );
  INV_X4 U117 ( .A(1'b1), .ZN(Output_MEMBus[78]) );
  INV_X4 U119 ( .A(1'b1), .ZN(Output_MEMBus[79]) );
  INV_X4 U121 ( .A(1'b1), .ZN(Output_MEMBus[80]) );
  INV_X4 U123 ( .A(1'b1), .ZN(Output_MEMBus[81]) );
  INV_X4 U125 ( .A(1'b1), .ZN(Output_MEMBus[82]) );
  INV_X4 U127 ( .A(1'b1), .ZN(Output_MEMBus[83]) );
  INV_X4 U129 ( .A(1'b1), .ZN(Output_MEMBus[84]) );
  INV_X4 U131 ( .A(1'b1), .ZN(Output_MEMBus[85]) );
  INV_X4 U133 ( .A(1'b1), .ZN(Output_MEMBus[86]) );
  INV_X4 U135 ( .A(1'b1), .ZN(Output_MEMBus[87]) );
  INV_X4 U137 ( .A(1'b1), .ZN(Output_MEMBus[88]) );
  INV_X4 U139 ( .A(1'b1), .ZN(Output_MEMBus[89]) );
  INV_X4 U141 ( .A(1'b1), .ZN(Output_MEMBus[90]) );
  INV_X4 U143 ( .A(1'b1), .ZN(Output_MEMBus[91]) );
  INV_X4 U145 ( .A(1'b1), .ZN(Output_MEMBus[92]) );
  INV_X4 U147 ( .A(1'b1), .ZN(Output_MEMBus[93]) );
  INV_X4 U149 ( .A(1'b1), .ZN(Output_MEMBus[94]) );
  INV_X4 U151 ( .A(1'b1), .ZN(Output_MEMBus[95]) );
  INV_X4 U153 ( .A(1'b1), .ZN(Output_MEMBus[96]) );
  INV_X4 U155 ( .A(1'b1), .ZN(Output_MEMBus[97]) );
  INV_X4 U157 ( .A(1'b1), .ZN(Output_MEMBus[98]) );
  INV_X4 U159 ( .A(1'b1), .ZN(Output_MEMBus[99]) );
  INV_X4 U161 ( .A(1'b1), .ZN(Output_MEMBus[100]) );
  INV_X4 U163 ( .A(1'b1), .ZN(Output_MEMBus[101]) );
  INV_X4 U165 ( .A(1'b1), .ZN(Output_MEMBus[102]) );
  INV_X4 U167 ( .A(1'b1), .ZN(Output_MEMBus[103]) );
  INV_X4 U169 ( .A(1'b1), .ZN(Output_MEMBus[104]) );
  INV_X4 U171 ( .A(1'b1), .ZN(Output_MEMBus[105]) );
  INV_X4 U173 ( .A(1'b1), .ZN(Output_MEMBus[106]) );
  INV_X4 U175 ( .A(1'b1), .ZN(Output_MEMBus[107]) );
  INV_X4 U177 ( .A(1'b1), .ZN(Output_MEMBus[108]) );
  INV_X4 U179 ( .A(1'b1), .ZN(Output_MEMBus[109]) );
  INV_X4 U181 ( .A(1'b1), .ZN(Output_MEMBus[110]) );
  INV_X4 U183 ( .A(1'b1), .ZN(Output_MEMBus[111]) );
  INV_X4 U185 ( .A(1'b1), .ZN(Output_MEMBus[112]) );
  INV_X4 U187 ( .A(1'b1), .ZN(Output_MEMBus[113]) );
  INV_X4 U189 ( .A(1'b1), .ZN(Output_MEMBus[114]) );
  INV_X4 U191 ( .A(1'b1), .ZN(Output_MEMBus[115]) );
  INV_X4 U193 ( .A(1'b1), .ZN(Output_MEMBus[116]) );
  INV_X4 U195 ( .A(1'b1), .ZN(Output_MEMBus[117]) );
  INV_X4 U197 ( .A(1'b1), .ZN(Output_MEMBus[118]) );
  INV_X4 U199 ( .A(1'b1), .ZN(Output_MEMBus[119]) );
  INV_X4 U201 ( .A(1'b1), .ZN(Output_MEMBus[120]) );
  INV_X4 U203 ( .A(1'b1), .ZN(Output_MEMBus[121]) );
  INV_X4 U205 ( .A(1'b1), .ZN(Output_MEMBus[122]) );
  INV_X4 U207 ( .A(1'b1), .ZN(Output_MEMBus[123]) );
  INV_X4 U209 ( .A(1'b1), .ZN(Output_MEMBus[124]) );
  INV_X4 U211 ( .A(1'b1), .ZN(Output_MEMBus[125]) );
  INV_X4 U213 ( .A(1'b1), .ZN(Output_MEMBus[126]) );
  INV_X4 U215 ( .A(1'b1), .ZN(Output_MEMBus[127]) );
  INV_X4 U217 ( .A(n218), .ZN(n217) );
  INV_X4 U218 ( .A(reset_n), .ZN(n218) );
endmodule


module input_top ( start, clock, rst_n, m1ReadBus, m2ReadBus, inputBaseOffset, 
        m1ReadAddr, m2ReadAddr, m2WriteAddr, m3WriteAddr, m2WriteBus, 
        m3WriteBus, m2WE, m3WE, done, cdf_valid, cdf_min );
  input [127:0] m1ReadBus;
  input [35:0] m2ReadBus;
  output [15:0] m1ReadAddr;
  output [15:0] m2ReadAddr;
  output [15:0] m2WriteAddr;
  output [15:0] m3WriteAddr;
  output [127:0] m2WriteBus;
  output [127:0] m3WriteBus;
  output [19:0] cdf_min;
  input start, clock, rst_n, inputBaseOffset;
  output m2WE, m3WE, done, cdf_valid;
  wire   n331, \U5/Z_0 , \U5/Z_1 , \U5/Z_2 , \U5/Z_3 , \U5/Z_4 , \U5/Z_5 ,
         \U5/Z_6 , \U5/Z_7 , \U5/Z_15 , \U5/DATA2_0 , \U5/DATA2_1 ,
         \U5/DATA2_2 , \U5/DATA2_3 , \U5/DATA2_4 , \U5/DATA2_5 , \U5/DATA2_6 ,
         \U5/DATA2_7 , \U5/DATA2_15 , \U5/DATA1_0 , \U5/DATA1_1 , \U5/DATA1_2 ,
         \U5/DATA1_3 , \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 , \U5/DATA1_7 ,
         \U5/DATA1_8 , \U5/DATA1_9 , \U5/DATA1_10 , \U5/DATA1_11 ,
         \U5/DATA1_12 , \U5/DATA1_13 , \U5/DATA1_14 , \U5/DATA1_15 , \U4/Z_0 ,
         \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 , \U4/Z_7 ,
         \U4/Z_8 , \U4/Z_9 , \U4/Z_10 , \U4/Z_11 , \U4/Z_12 , \U4/Z_13 ,
         \U4/Z_14 , \U4/Z_15 , \U4/Z_16 , \U4/Z_17 , \U4/Z_18 , \U4/Z_19 ,
         \U4/DATA2_0 , \U4/DATA2_1 , \U4/DATA2_2 , \U4/DATA2_3 , \U4/DATA2_4 ,
         \U4/DATA2_5 , \U4/DATA2_6 , \U4/DATA2_7 , \U4/DATA2_8 , \U4/DATA2_9 ,
         \U4/DATA2_10 , \U4/DATA2_11 , \U4/DATA2_12 , \U4/DATA2_13 ,
         \U4/DATA2_14 , \U4/DATA2_15 , \U4/DATA2_16 , \U4/DATA2_17 ,
         \U4/DATA2_18 , \U4/DATA2_19 , \U4/DATA2_20 , \U4/DATA2_21 ,
         \U4/DATA2_22 , \U4/DATA2_23 , \U4/DATA2_24 , \U4/DATA2_25 ,
         \U4/DATA2_26 , \U4/DATA2_27 , \U4/DATA2_28 , \U4/DATA2_29 ,
         \U4/DATA2_30 , \U4/DATA2_31 , \U4/DATA2_32 , \U4/DATA2_33 ,
         \U4/DATA2_34 , \U4/DATA2_35 , \U4/DATA1_0 , \U4/DATA1_1 ,
         \U4/DATA1_2 , \U4/DATA1_3 , \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 ,
         \U4/DATA1_7 , \U4/DATA1_8 , \U4/DATA1_9 , \U4/DATA1_10 ,
         \U4/DATA1_11 , \U4/DATA1_12 , \U4/DATA1_13 , \U4/DATA1_14 ,
         \U4/DATA1_15 , \U4/DATA1_16 , \U4/DATA1_17 , \U4/DATA1_18 ,
         \U4/DATA1_19 , \U3/Z_0 , \U3/Z_1 , \U3/Z_2 , \U3/Z_3 , \U3/Z_4 ,
         \U3/Z_5 , \U3/Z_6 , \U3/Z_7 , \U3/Z_15 , \U3/DATA2_0 , \U3/DATA2_1 ,
         \U3/DATA2_2 , \U3/DATA2_3 , \U3/DATA2_4 , \U3/DATA2_5 , \U3/DATA2_6 ,
         \U3/DATA2_7 , \U3/DATA2_15 , \U3/DATA1_0 , \U3/DATA1_1 , \U3/DATA1_2 ,
         \U3/DATA1_3 , \U3/DATA1_4 , \U3/DATA1_5 , \U3/DATA1_6 , \U3/DATA1_7 ,
         \U3/DATA1_8 , \U3/DATA1_9 , \U3/DATA1_10 , \U3/DATA1_11 ,
         \U3/DATA1_12 , \U3/DATA1_13 , \U3/DATA1_14 , \U3/DATA1_15 , \U2/Z_0 ,
         \U2/DATA2_0 , \U2/DATA1_0 , n165, n166, n167, n168, n169, n170, n171,
         n177, n178, n189, n200, n211, n222, n233, n244, n255, n266, n267,
         n268, n269, n270, n271, n272, n273, n282, n293, n304, n305, n306,
         n309, n310, n311, n312, n313, n314, n315, n321, n322, n323, n1158,
         n1159, n1160, n1161;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213;
  assign m2WriteAddr[0] = \U5/Z_0 ;
  assign m2WriteAddr[1] = \U5/Z_1 ;
  assign m2WriteAddr[2] = \U5/Z_2 ;
  assign m2WriteAddr[3] = \U5/Z_3 ;
  assign m2WriteAddr[4] = \U5/Z_4 ;
  assign m2WriteAddr[5] = \U5/Z_5 ;
  assign m2WriteAddr[6] = \U5/Z_6 ;
  assign m2WriteAddr[7] = \U5/Z_7 ;
  assign m2WriteAddr[15] = \U5/Z_15 ;
  assign m2WriteBus[0] = \U4/Z_0 ;
  assign m2WriteBus[1] = \U4/Z_1 ;
  assign m2WriteBus[2] = \U4/Z_2 ;
  assign m2WriteBus[3] = \U4/Z_3 ;
  assign m2WriteBus[4] = \U4/Z_4 ;
  assign m2WriteBus[5] = \U4/Z_5 ;
  assign m2WriteBus[6] = \U4/Z_6 ;
  assign m2WriteBus[7] = \U4/Z_7 ;
  assign m2WriteBus[8] = \U4/Z_8 ;
  assign m2WriteBus[9] = \U4/Z_9 ;
  assign m2WriteBus[10] = \U4/Z_10 ;
  assign m2WriteBus[11] = \U4/Z_11 ;
  assign m2WriteBus[12] = \U4/Z_12 ;
  assign m2WriteBus[13] = \U4/Z_13 ;
  assign m2WriteBus[14] = \U4/Z_14 ;
  assign m2WriteBus[15] = \U4/Z_15 ;
  assign m2WriteBus[16] = \U4/Z_16 ;
  assign m2WriteBus[17] = \U4/Z_17 ;
  assign m2WriteBus[18] = \U4/Z_18 ;
  assign m2WriteBus[19] = \U4/Z_19 ;
  assign m2ReadAddr[0] = \U3/Z_0 ;
  assign m2ReadAddr[1] = \U3/Z_1 ;
  assign m2ReadAddr[2] = \U3/Z_2 ;
  assign m2ReadAddr[3] = \U3/Z_3 ;
  assign m2ReadAddr[4] = \U3/Z_4 ;
  assign m2ReadAddr[5] = \U3/Z_5 ;
  assign m2ReadAddr[6] = \U3/Z_6 ;
  assign m2ReadAddr[7] = \U3/Z_7 ;
  assign m2ReadAddr[15] = \U3/Z_15 ;
  assign m2WE = \U2/Z_0 ;

  INV_X4 U5 ( .A(n165), .ZN(\U5/Z_7 ) );
  INV_X4 U7 ( .A(n166), .ZN(\U5/Z_6 ) );
  INV_X4 U9 ( .A(n167), .ZN(\U5/Z_5 ) );
  INV_X4 U11 ( .A(n168), .ZN(\U5/Z_4 ) );
  INV_X4 U13 ( .A(n169), .ZN(\U5/Z_3 ) );
  INV_X4 U15 ( .A(n170), .ZN(\U5/Z_2 ) );
  INV_X4 U17 ( .A(n171), .ZN(\U5/Z_15 ) );
  INV_X4 U29 ( .A(n177), .ZN(\U5/Z_1 ) );
  INV_X4 U31 ( .A(n178), .ZN(\U5/Z_0 ) );
  INV_X4 U53 ( .A(n189), .ZN(\U4/Z_9 ) );
  INV_X4 U75 ( .A(n200), .ZN(\U4/Z_8 ) );
  INV_X4 U97 ( .A(n211), .ZN(\U4/Z_7 ) );
  INV_X4 U119 ( .A(n222), .ZN(\U4/Z_6 ) );
  INV_X4 U141 ( .A(n233), .ZN(\U4/Z_5 ) );
  INV_X4 U163 ( .A(n244), .ZN(\U4/Z_4 ) );
  INV_X4 U185 ( .A(n255), .ZN(\U4/Z_3 ) );
  INV_X4 U207 ( .A(n266), .ZN(\U4/Z_2 ) );
  INV_X4 U209 ( .A(n267), .ZN(\U4/Z_19 ) );
  INV_X4 U211 ( .A(n268), .ZN(\U4/Z_18 ) );
  INV_X4 U213 ( .A(n269), .ZN(\U4/Z_17 ) );
  INV_X4 U215 ( .A(n270), .ZN(\U4/Z_16 ) );
  INV_X4 U217 ( .A(n271), .ZN(\U4/Z_15 ) );
  INV_X4 U219 ( .A(n272), .ZN(\U4/Z_14 ) );
  INV_X4 U221 ( .A(n273), .ZN(\U4/Z_13 ) );
  INV_X4 U239 ( .A(n282), .ZN(\U4/Z_12 ) );
  INV_X4 U261 ( .A(n293), .ZN(\U4/Z_11 ) );
  INV_X4 U283 ( .A(n304), .ZN(\U4/Z_10 ) );
  INV_X4 U285 ( .A(n305), .ZN(\U4/Z_1 ) );
  INV_X4 U287 ( .A(n306), .ZN(\U4/Z_0 ) );
  INV_X4 U293 ( .A(n309), .ZN(\U3/Z_7 ) );
  INV_X4 U295 ( .A(n310), .ZN(\U3/Z_6 ) );
  INV_X4 U297 ( .A(n311), .ZN(\U3/Z_5 ) );
  INV_X4 U299 ( .A(n312), .ZN(\U3/Z_4 ) );
  INV_X4 U301 ( .A(n313), .ZN(\U3/Z_3 ) );
  INV_X4 U303 ( .A(n314), .ZN(\U3/Z_2 ) );
  INV_X4 U305 ( .A(n315), .ZN(\U3/Z_15 ) );
  INV_X4 U317 ( .A(n321), .ZN(\U3/Z_1 ) );
  INV_X4 U319 ( .A(n322), .ZN(\U3/Z_0 ) );
  INV_X4 U321 ( .A(n323), .ZN(\U2/Z_0 ) );
  input_pipeline input_dut ( .start(start), .clock(clock), .rst_n(n1160), 
        .m1ReadBus(m1ReadBus), .m2ReadBus(m2ReadBus), .inputBaseOffset(
        inputBaseOffset), .m1ReadAddr(m1ReadAddr), .m2ReadAddr({\U3/DATA2_15 , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, \U3/DATA2_7 , \U3/DATA2_6 , \U3/DATA2_5 , 
        \U3/DATA2_4 , \U3/DATA2_3 , \U3/DATA2_2 , \U3/DATA2_1 , \U3/DATA2_0 }), 
        .m2WriteAddr({\U5/DATA2_15 , SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, \U5/DATA2_7 , 
        \U5/DATA2_6 , \U5/DATA2_5 , \U5/DATA2_4 , \U5/DATA2_3 , \U5/DATA2_2 , 
        \U5/DATA2_1 , \U5/DATA2_0 }), .m3WriteAddr(m3WriteAddr), .m2WriteBus({
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, \U4/DATA2_35 , 
        \U4/DATA2_34 , \U4/DATA2_33 , \U4/DATA2_32 , \U4/DATA2_31 , 
        \U4/DATA2_30 , \U4/DATA2_29 , \U4/DATA2_28 , \U4/DATA2_27 , 
        \U4/DATA2_26 , \U4/DATA2_25 , \U4/DATA2_24 , \U4/DATA2_23 , 
        \U4/DATA2_22 , \U4/DATA2_21 , \U4/DATA2_20 , \U4/DATA2_19 , 
        \U4/DATA2_18 , \U4/DATA2_17 , \U4/DATA2_16 , \U4/DATA2_15 , 
        \U4/DATA2_14 , \U4/DATA2_13 , \U4/DATA2_12 , \U4/DATA2_11 , 
        \U4/DATA2_10 , \U4/DATA2_9 , \U4/DATA2_8 , \U4/DATA2_7 , \U4/DATA2_6 , 
        \U4/DATA2_5 , \U4/DATA2_4 , \U4/DATA2_3 , \U4/DATA2_2 , \U4/DATA2_1 , 
        \U4/DATA2_0 }), .m3WriteBus(m3WriteBus), .m2WE(\U2/DATA2_0 ), .m3WE(
        m3WE), .input_done(n331) );
  Cdf_top CDF_dut ( .clock(clock), .reset_n(n1160), .start(n1158), 
        .SP_ReadBus(m2ReadBus), .SP_ReadAddress({\U3/DATA1_15 , \U3/DATA1_14 , 
        \U3/DATA1_13 , \U3/DATA1_12 , \U3/DATA1_11 , \U3/DATA1_10 , 
        \U3/DATA1_9 , \U3/DATA1_8 , \U3/DATA1_7 , \U3/DATA1_6 , \U3/DATA1_5 , 
        \U3/DATA1_4 , \U3/DATA1_3 , \U3/DATA1_2 , \U3/DATA1_1 , \U3/DATA1_0 }), 
        .WriteEnable(\U2/DATA1_0 ), .Output_MEMBus({SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, 
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, 
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        SYNOPSYS_UNCONNECTED__151, SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, 
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, 
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, 
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, SYNOPSYS_UNCONNECTED__186, 
        SYNOPSYS_UNCONNECTED__187, SYNOPSYS_UNCONNECTED__188, 
        SYNOPSYS_UNCONNECTED__189, SYNOPSYS_UNCONNECTED__190, 
        SYNOPSYS_UNCONNECTED__191, SYNOPSYS_UNCONNECTED__192, 
        SYNOPSYS_UNCONNECTED__193, SYNOPSYS_UNCONNECTED__194, 
        SYNOPSYS_UNCONNECTED__195, SYNOPSYS_UNCONNECTED__196, 
        SYNOPSYS_UNCONNECTED__197, SYNOPSYS_UNCONNECTED__198, 
        SYNOPSYS_UNCONNECTED__199, SYNOPSYS_UNCONNECTED__200, 
        SYNOPSYS_UNCONNECTED__201, SYNOPSYS_UNCONNECTED__202, 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, 
        SYNOPSYS_UNCONNECTED__207, SYNOPSYS_UNCONNECTED__208, 
        SYNOPSYS_UNCONNECTED__209, SYNOPSYS_UNCONNECTED__210, 
        SYNOPSYS_UNCONNECTED__211, SYNOPSYS_UNCONNECTED__212, 
        SYNOPSYS_UNCONNECTED__213, \U4/DATA1_19 , \U4/DATA1_18 , \U4/DATA1_17 , 
        \U4/DATA1_16 , \U4/DATA1_15 , \U4/DATA1_14 , \U4/DATA1_13 , 
        \U4/DATA1_12 , \U4/DATA1_11 , \U4/DATA1_10 , \U4/DATA1_9 , 
        \U4/DATA1_8 , \U4/DATA1_7 , \U4/DATA1_6 , \U4/DATA1_5 , \U4/DATA1_4 , 
        \U4/DATA1_3 , \U4/DATA1_2 , \U4/DATA1_1 , \U4/DATA1_0 }), 
        .Output_MEMAddress({\U5/DATA1_15 , \U5/DATA1_14 , \U5/DATA1_13 , 
        \U5/DATA1_12 , \U5/DATA1_11 , \U5/DATA1_10 , \U5/DATA1_9 , 
        \U5/DATA1_8 , \U5/DATA1_7 , \U5/DATA1_6 , \U5/DATA1_5 , \U5/DATA1_4 , 
        \U5/DATA1_3 , \U5/DATA1_2 , \U5/DATA1_1 , \U5/DATA1_0 }), .Cdf_Min(
        cdf_min), .done(done), .input_base_offset(inputBaseOffset), 
        .cdf_valid(cdf_valid) );
  INV_X4 U1 ( .A(1'b1), .ZN(m2WriteBus[36]) );
  INV_X4 U3 ( .A(1'b1), .ZN(m2WriteBus[37]) );
  INV_X4 U6 ( .A(1'b1), .ZN(m2WriteBus[38]) );
  INV_X4 U10 ( .A(1'b1), .ZN(m2WriteBus[39]) );
  INV_X4 U14 ( .A(1'b1), .ZN(m2WriteBus[40]) );
  INV_X4 U18 ( .A(1'b1), .ZN(m2WriteBus[41]) );
  INV_X4 U20 ( .A(1'b1), .ZN(m2WriteBus[42]) );
  INV_X4 U22 ( .A(1'b1), .ZN(m2WriteBus[43]) );
  INV_X4 U24 ( .A(1'b1), .ZN(m2WriteBus[44]) );
  INV_X4 U26 ( .A(1'b1), .ZN(m2WriteBus[45]) );
  INV_X4 U28 ( .A(1'b1), .ZN(m2WriteBus[46]) );
  INV_X4 U32 ( .A(1'b1), .ZN(m2WriteBus[47]) );
  INV_X4 U34 ( .A(1'b1), .ZN(m2WriteBus[48]) );
  INV_X4 U36 ( .A(1'b1), .ZN(m2WriteBus[49]) );
  INV_X4 U38 ( .A(1'b1), .ZN(m2WriteBus[50]) );
  INV_X4 U40 ( .A(1'b1), .ZN(m2WriteBus[51]) );
  INV_X4 U42 ( .A(1'b1), .ZN(m2WriteBus[52]) );
  INV_X4 U44 ( .A(1'b1), .ZN(m2WriteBus[53]) );
  INV_X4 U46 ( .A(1'b1), .ZN(m2WriteBus[54]) );
  INV_X4 U48 ( .A(1'b1), .ZN(m2WriteBus[55]) );
  INV_X4 U50 ( .A(1'b1), .ZN(m2WriteBus[56]) );
  INV_X4 U52 ( .A(1'b1), .ZN(m2WriteBus[57]) );
  INV_X4 U55 ( .A(1'b1), .ZN(m2WriteBus[58]) );
  INV_X4 U57 ( .A(1'b1), .ZN(m2WriteBus[59]) );
  INV_X4 U59 ( .A(1'b1), .ZN(m2WriteBus[60]) );
  INV_X4 U61 ( .A(1'b1), .ZN(m2WriteBus[61]) );
  INV_X4 U63 ( .A(1'b1), .ZN(m2WriteBus[62]) );
  INV_X4 U65 ( .A(1'b1), .ZN(m2WriteBus[63]) );
  INV_X4 U67 ( .A(1'b1), .ZN(m2WriteBus[64]) );
  INV_X4 U69 ( .A(1'b1), .ZN(m2WriteBus[65]) );
  INV_X4 U71 ( .A(1'b1), .ZN(m2WriteBus[66]) );
  INV_X4 U73 ( .A(1'b1), .ZN(m2WriteBus[67]) );
  INV_X4 U76 ( .A(1'b1), .ZN(m2WriteBus[68]) );
  INV_X4 U78 ( .A(1'b1), .ZN(m2WriteBus[69]) );
  INV_X4 U80 ( .A(1'b1), .ZN(m2WriteBus[70]) );
  INV_X4 U82 ( .A(1'b1), .ZN(m2WriteBus[71]) );
  INV_X4 U84 ( .A(1'b1), .ZN(m2WriteBus[72]) );
  INV_X4 U86 ( .A(1'b1), .ZN(m2WriteBus[73]) );
  INV_X4 U88 ( .A(1'b1), .ZN(m2WriteBus[74]) );
  INV_X4 U90 ( .A(1'b1), .ZN(m2WriteBus[75]) );
  INV_X4 U92 ( .A(1'b1), .ZN(m2WriteBus[76]) );
  INV_X4 U94 ( .A(1'b1), .ZN(m2WriteBus[77]) );
  INV_X4 U96 ( .A(1'b1), .ZN(m2WriteBus[78]) );
  INV_X4 U99 ( .A(1'b1), .ZN(m2WriteBus[79]) );
  INV_X4 U101 ( .A(1'b1), .ZN(m2WriteBus[80]) );
  INV_X4 U103 ( .A(1'b1), .ZN(m2WriteBus[81]) );
  INV_X4 U105 ( .A(1'b1), .ZN(m2WriteBus[82]) );
  INV_X4 U107 ( .A(1'b1), .ZN(m2WriteBus[83]) );
  INV_X4 U109 ( .A(1'b1), .ZN(m2WriteBus[84]) );
  INV_X4 U111 ( .A(1'b1), .ZN(m2WriteBus[85]) );
  INV_X4 U113 ( .A(1'b1), .ZN(m2WriteBus[86]) );
  INV_X4 U115 ( .A(1'b1), .ZN(m2WriteBus[87]) );
  INV_X4 U117 ( .A(1'b1), .ZN(m2WriteBus[88]) );
  INV_X4 U120 ( .A(1'b1), .ZN(m2WriteBus[89]) );
  INV_X4 U122 ( .A(1'b1), .ZN(m2WriteBus[90]) );
  INV_X4 U124 ( .A(1'b1), .ZN(m2WriteBus[91]) );
  INV_X4 U126 ( .A(1'b1), .ZN(m2WriteBus[92]) );
  INV_X4 U128 ( .A(1'b1), .ZN(m2WriteBus[93]) );
  INV_X4 U130 ( .A(1'b1), .ZN(m2WriteBus[94]) );
  INV_X4 U132 ( .A(1'b1), .ZN(m2WriteBus[95]) );
  INV_X4 U134 ( .A(1'b1), .ZN(m2WriteBus[96]) );
  INV_X4 U136 ( .A(1'b1), .ZN(m2WriteBus[97]) );
  INV_X4 U138 ( .A(1'b1), .ZN(m2WriteBus[98]) );
  INV_X4 U140 ( .A(1'b1), .ZN(m2WriteBus[99]) );
  INV_X4 U143 ( .A(1'b1), .ZN(m2WriteBus[100]) );
  INV_X4 U145 ( .A(1'b1), .ZN(m2WriteBus[101]) );
  INV_X4 U147 ( .A(1'b1), .ZN(m2WriteBus[102]) );
  INV_X4 U149 ( .A(1'b1), .ZN(m2WriteBus[103]) );
  INV_X4 U151 ( .A(1'b1), .ZN(m2WriteBus[104]) );
  INV_X4 U153 ( .A(1'b1), .ZN(m2WriteBus[105]) );
  INV_X4 U155 ( .A(1'b1), .ZN(m2WriteBus[106]) );
  INV_X4 U157 ( .A(1'b1), .ZN(m2WriteBus[107]) );
  INV_X4 U159 ( .A(1'b1), .ZN(m2WriteBus[108]) );
  INV_X4 U161 ( .A(1'b1), .ZN(m2WriteBus[109]) );
  INV_X4 U164 ( .A(1'b1), .ZN(m2WriteBus[110]) );
  INV_X4 U166 ( .A(1'b1), .ZN(m2WriteBus[111]) );
  INV_X4 U168 ( .A(1'b1), .ZN(m2WriteBus[112]) );
  INV_X4 U170 ( .A(1'b1), .ZN(m2WriteBus[113]) );
  INV_X4 U172 ( .A(1'b1), .ZN(m2WriteBus[114]) );
  INV_X4 U174 ( .A(1'b1), .ZN(m2WriteBus[115]) );
  INV_X4 U176 ( .A(1'b1), .ZN(m2WriteBus[116]) );
  INV_X4 U178 ( .A(1'b1), .ZN(m2WriteBus[117]) );
  INV_X4 U180 ( .A(1'b1), .ZN(m2WriteBus[118]) );
  INV_X4 U182 ( .A(1'b1), .ZN(m2WriteBus[119]) );
  INV_X4 U184 ( .A(1'b1), .ZN(m2WriteBus[120]) );
  INV_X4 U187 ( .A(1'b1), .ZN(m2WriteBus[121]) );
  INV_X4 U189 ( .A(1'b1), .ZN(m2WriteBus[122]) );
  INV_X4 U191 ( .A(1'b1), .ZN(m2WriteBus[123]) );
  INV_X4 U193 ( .A(1'b1), .ZN(m2WriteBus[124]) );
  INV_X4 U195 ( .A(1'b1), .ZN(m2WriteBus[125]) );
  INV_X4 U197 ( .A(1'b1), .ZN(m2WriteBus[126]) );
  INV_X4 U199 ( .A(1'b1), .ZN(m2WriteBus[127]) );
  AND2_X4 U201 ( .A1(\U4/DATA2_20 ), .A2(n1159), .ZN(m2WriteBus[20]) );
  AND2_X4 U202 ( .A1(\U4/DATA2_21 ), .A2(n1159), .ZN(m2WriteBus[21]) );
  AND2_X4 U203 ( .A1(\U4/DATA2_22 ), .A2(n1159), .ZN(m2WriteBus[22]) );
  AND2_X4 U204 ( .A1(\U4/DATA2_23 ), .A2(n1159), .ZN(m2WriteBus[23]) );
  AND2_X4 U205 ( .A1(\U4/DATA2_24 ), .A2(n1159), .ZN(m2WriteBus[24]) );
  AND2_X4 U206 ( .A1(\U4/DATA2_25 ), .A2(n1159), .ZN(m2WriteBus[25]) );
  AND2_X4 U208 ( .A1(\U4/DATA2_26 ), .A2(n1159), .ZN(m2WriteBus[26]) );
  AND2_X4 U210 ( .A1(\U4/DATA2_27 ), .A2(n1159), .ZN(m2WriteBus[27]) );
  AND2_X4 U212 ( .A1(\U4/DATA2_28 ), .A2(n1159), .ZN(m2WriteBus[28]) );
  AND2_X4 U214 ( .A1(\U4/DATA2_29 ), .A2(n1159), .ZN(m2WriteBus[29]) );
  AND2_X4 U216 ( .A1(\U4/DATA2_30 ), .A2(n1159), .ZN(m2WriteBus[30]) );
  AND2_X4 U218 ( .A1(\U4/DATA2_31 ), .A2(n1159), .ZN(m2WriteBus[31]) );
  AND2_X4 U220 ( .A1(\U4/DATA2_32 ), .A2(n1159), .ZN(m2WriteBus[32]) );
  AND2_X4 U222 ( .A1(\U4/DATA2_33 ), .A2(n1159), .ZN(m2WriteBus[33]) );
  AND2_X4 U223 ( .A1(\U4/DATA2_34 ), .A2(n1159), .ZN(m2WriteBus[34]) );
  AND2_X4 U224 ( .A1(\U4/DATA2_35 ), .A2(n1159), .ZN(m2WriteBus[35]) );
  AND2_X4 U225 ( .A1(\U5/DATA1_8 ), .A2(n331), .ZN(m2WriteAddr[8]) );
  AND2_X4 U226 ( .A1(\U5/DATA1_10 ), .A2(n331), .ZN(m2WriteAddr[10]) );
  AND2_X4 U227 ( .A1(\U5/DATA1_11 ), .A2(n331), .ZN(m2WriteAddr[11]) );
  AND2_X4 U228 ( .A1(\U5/DATA1_12 ), .A2(n331), .ZN(m2WriteAddr[12]) );
  AND2_X4 U229 ( .A1(\U5/DATA1_13 ), .A2(n331), .ZN(m2WriteAddr[13]) );
  AND2_X4 U230 ( .A1(\U5/DATA1_14 ), .A2(n331), .ZN(m2WriteAddr[14]) );
  AND2_X4 U231 ( .A1(\U3/DATA1_14 ), .A2(n331), .ZN(m2ReadAddr[14]) );
  AND2_X4 U232 ( .A1(n1158), .A2(\U5/DATA1_9 ), .ZN(m2WriteAddr[9]) );
  AND2_X4 U233 ( .A1(\U3/DATA1_12 ), .A2(n331), .ZN(m2ReadAddr[12]) );
  AND2_X4 U234 ( .A1(\U3/DATA1_13 ), .A2(n331), .ZN(m2ReadAddr[13]) );
  AND2_X4 U235 ( .A1(\U3/DATA1_8 ), .A2(n331), .ZN(m2ReadAddr[8]) );
  AND2_X4 U236 ( .A1(\U3/DATA1_9 ), .A2(n331), .ZN(m2ReadAddr[9]) );
  AND2_X4 U237 ( .A1(\U3/DATA1_10 ), .A2(n331), .ZN(m2ReadAddr[10]) );
  AND2_X4 U238 ( .A1(\U3/DATA1_11 ), .A2(n331), .ZN(m2ReadAddr[11]) );
  INV_X4 U240 ( .A(n1159), .ZN(n1158) );
  INV_X4 U241 ( .A(n1161), .ZN(n1160) );
  INV_X4 U242 ( .A(rst_n), .ZN(n1161) );
  AOI22_X2 U243 ( .A1(\U4/DATA1_0 ), .A2(n1158), .B1(\U4/DATA2_0 ), .B2(n1159), 
        .ZN(n306) );
  AOI22_X2 U244 ( .A1(\U4/DATA1_1 ), .A2(n1158), .B1(\U4/DATA2_1 ), .B2(n1159), 
        .ZN(n305) );
  AOI22_X2 U245 ( .A1(\U4/DATA1_10 ), .A2(n1158), .B1(\U4/DATA2_10 ), .B2(
        n1159), .ZN(n304) );
  AOI22_X2 U246 ( .A1(\U4/DATA1_11 ), .A2(n1158), .B1(\U4/DATA2_11 ), .B2(
        n1159), .ZN(n293) );
  AOI22_X2 U247 ( .A1(\U4/DATA1_12 ), .A2(n1158), .B1(\U4/DATA2_12 ), .B2(
        n1159), .ZN(n282) );
  AOI22_X2 U248 ( .A1(\U4/DATA1_13 ), .A2(n1158), .B1(\U4/DATA2_13 ), .B2(
        n1159), .ZN(n273) );
  AOI22_X2 U249 ( .A1(\U4/DATA1_14 ), .A2(n1158), .B1(\U4/DATA2_14 ), .B2(
        n1159), .ZN(n272) );
  AOI22_X2 U250 ( .A1(\U4/DATA1_15 ), .A2(n1158), .B1(\U4/DATA2_15 ), .B2(
        n1159), .ZN(n271) );
  AOI22_X2 U251 ( .A1(\U4/DATA1_16 ), .A2(n1158), .B1(\U4/DATA2_16 ), .B2(
        n1159), .ZN(n270) );
  AOI22_X2 U252 ( .A1(\U4/DATA1_17 ), .A2(n331), .B1(\U4/DATA2_17 ), .B2(n1159), .ZN(n269) );
  AOI22_X2 U253 ( .A1(\U4/DATA1_18 ), .A2(n331), .B1(\U4/DATA2_18 ), .B2(n1159), .ZN(n268) );
  AOI22_X2 U254 ( .A1(\U4/DATA1_2 ), .A2(n1158), .B1(\U4/DATA2_2 ), .B2(n1159), 
        .ZN(n266) );
  AOI22_X2 U255 ( .A1(\U4/DATA1_3 ), .A2(n1158), .B1(\U4/DATA2_3 ), .B2(n1159), 
        .ZN(n255) );
  AOI22_X2 U256 ( .A1(\U4/DATA1_4 ), .A2(n1158), .B1(\U4/DATA2_4 ), .B2(n1159), 
        .ZN(n244) );
  AOI22_X2 U257 ( .A1(\U4/DATA1_5 ), .A2(n331), .B1(\U4/DATA2_5 ), .B2(n1159), 
        .ZN(n233) );
  AOI22_X2 U258 ( .A1(\U4/DATA1_6 ), .A2(n1158), .B1(\U4/DATA2_6 ), .B2(n1159), 
        .ZN(n222) );
  AOI22_X2 U259 ( .A1(\U4/DATA1_7 ), .A2(n331), .B1(\U4/DATA2_7 ), .B2(n1159), 
        .ZN(n211) );
  AOI22_X2 U260 ( .A1(\U4/DATA1_8 ), .A2(n1158), .B1(\U4/DATA2_8 ), .B2(n1159), 
        .ZN(n200) );
  AOI22_X2 U262 ( .A1(\U4/DATA1_9 ), .A2(n331), .B1(\U4/DATA2_9 ), .B2(n1159), 
        .ZN(n189) );
  AOI22_X2 U263 ( .A1(\U4/DATA1_19 ), .A2(n1158), .B1(\U4/DATA2_19 ), .B2(
        n1159), .ZN(n267) );
  INV_X4 U264 ( .A(n331), .ZN(n1159) );
  AOI22_X2 U265 ( .A1(\U5/DATA1_4 ), .A2(n331), .B1(\U5/DATA2_4 ), .B2(n1159), 
        .ZN(n168) );
  AOI22_X2 U266 ( .A1(\U5/DATA1_5 ), .A2(n1158), .B1(\U5/DATA2_5 ), .B2(n1159), 
        .ZN(n167) );
  AOI22_X2 U267 ( .A1(\U5/DATA1_6 ), .A2(n331), .B1(\U5/DATA2_6 ), .B2(n1159), 
        .ZN(n166) );
  AOI22_X2 U268 ( .A1(\U5/DATA1_7 ), .A2(n1158), .B1(\U5/DATA2_7 ), .B2(n1159), 
        .ZN(n165) );
  AOI22_X2 U269 ( .A1(\U2/DATA1_0 ), .A2(n331), .B1(\U2/DATA2_0 ), .B2(n1159), 
        .ZN(n323) );
  AOI22_X1 U270 ( .A1(\U3/DATA1_0 ), .A2(n331), .B1(\U3/DATA2_0 ), .B2(n1159), 
        .ZN(n322) );
  AOI22_X1 U271 ( .A1(\U3/DATA1_1 ), .A2(n331), .B1(\U3/DATA2_1 ), .B2(n1159), 
        .ZN(n321) );
  AOI22_X2 U272 ( .A1(\U3/DATA1_3 ), .A2(n1158), .B1(\U3/DATA2_3 ), .B2(n1159), 
        .ZN(n313) );
  AOI22_X2 U273 ( .A1(\U3/DATA1_4 ), .A2(n331), .B1(\U3/DATA2_4 ), .B2(n1159), 
        .ZN(n312) );
  AOI22_X2 U274 ( .A1(\U3/DATA1_5 ), .A2(n331), .B1(\U3/DATA2_5 ), .B2(n1159), 
        .ZN(n311) );
  AOI22_X2 U275 ( .A1(\U3/DATA1_6 ), .A2(n331), .B1(\U3/DATA2_6 ), .B2(n1159), 
        .ZN(n310) );
  AOI22_X2 U276 ( .A1(\U3/DATA1_7 ), .A2(n331), .B1(\U3/DATA2_7 ), .B2(n1159), 
        .ZN(n309) );
  AOI22_X2 U277 ( .A1(\U5/DATA1_0 ), .A2(n331), .B1(\U5/DATA2_0 ), .B2(n1159), 
        .ZN(n178) );
  AOI22_X2 U278 ( .A1(\U5/DATA1_1 ), .A2(n1158), .B1(\U5/DATA2_1 ), .B2(n1159), 
        .ZN(n177) );
  AOI22_X2 U279 ( .A1(\U5/DATA1_2 ), .A2(n331), .B1(\U5/DATA2_2 ), .B2(n1159), 
        .ZN(n170) );
  AOI22_X2 U280 ( .A1(\U5/DATA1_3 ), .A2(n1158), .B1(\U5/DATA2_3 ), .B2(n1159), 
        .ZN(n169) );
  AOI22_X2 U281 ( .A1(\U5/DATA1_15 ), .A2(n331), .B1(\U5/DATA2_15 ), .B2(n1159), .ZN(n171) );
  AOI22_X2 U282 ( .A1(\U3/DATA1_2 ), .A2(n331), .B1(\U3/DATA2_2 ), .B2(n1159), 
        .ZN(n314) );
  AOI22_X2 U284 ( .A1(\U3/DATA1_15 ), .A2(n1158), .B1(\U3/DATA2_15 ), .B2(
        n1159), .ZN(n315) );
endmodule


module Top ( clock, reset_n, start, M1_ReadBus1, M1_ReadAddress1, M2_ReadBus1, 
        M2_ReadBus2, M2_ReadAddress1, M2_ReadAddress2, M2_WriteBus, 
        M2_WriteAddress, M2_WriteEnable, M3_ReadBus1, M3_ReadAddress1, 
        M3_WriteBus, M3_WriteAddress, M3_WriteEnable, M4_WriteBus, 
        M4_WriteAddress, M4_WriteEnable );
  input [127:0] M1_ReadBus1;
  output [15:0] M1_ReadAddress1;
  input [35:0] M2_ReadBus1;
  input [19:0] M2_ReadBus2;
  output [15:0] M2_ReadAddress1;
  output [15:0] M2_ReadAddress2;
  output [127:0] M2_WriteBus;
  output [15:0] M2_WriteAddress;
  input [127:0] M3_ReadBus1;
  output [15:0] M3_ReadAddress1;
  output [127:0] M3_WriteBus;
  output [15:0] M3_WriteAddress;
  output [127:0] M4_WriteBus;
  output [15:0] M4_WriteAddress;
  input clock, reset_n, start;
  output M2_WriteEnable, M3_WriteEnable, M4_WriteEnable;
  wire   input_base_offset, output_base_offset, output_start, input_start,
         output_done, input_done, cdf_valid, n200, n201;
  wire   [19:0] cdf_min;
  wire   [19:0] cdf_min_out;
  wire   [19:0] divisor;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98;

  Output_top dut_output_top ( .clock(clock), .reset_n(n200), .start(
        output_start), .CdfMin(cdf_min_out), .divisor(divisor), .M2SP_ReadBus(
        M2_ReadBus2), .M2SP_ReadAddress({M2_ReadAddress2[15], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, M2_ReadAddress2[7:0]}), .M3SP_ReadBus(
        M3_ReadBus1), .M3SP_ReadAddress(M3_ReadAddress1), .WriteEnable(
        M4_WriteEnable), .Output_MEMBus(M4_WriteBus), .Output_MEMAddress(
        M4_WriteAddress), .done(output_done), .output_base_offset(
        output_base_offset) );
  Controllor dut_Controller ( .clock(clock), .reset_n(n200), .start(start), 
        .output_start(output_start), .input_start(input_start), .input_done(
        input_done), .output_done(output_done), .Cdf_Min(cdf_min), 
        .Cdf_Min_Out(cdf_min_out), .Divisor(divisor), .output_base_offset(
        output_base_offset), .input_base_offset(input_base_offset), 
        .cdf_valid(cdf_valid) );
  input_top top_dut ( .start(input_start), .clock(clock), .rst_n(n200), 
        .m1ReadBus(M1_ReadBus1), .m2ReadBus(M2_ReadBus1), .inputBaseOffset(
        input_base_offset), .m1ReadAddr(M1_ReadAddress1), .m2ReadAddr(
        M2_ReadAddress1), .m2WriteAddr(M2_WriteAddress), .m3WriteAddr(
        M3_WriteAddress), .m2WriteBus({SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, M2_WriteBus[35:0]}), .m3WriteBus(M3_WriteBus), .m2WE(M2_WriteEnable), .m3WE(M3_WriteEnable), .done(input_done), .cdf_valid(
        cdf_valid), .cdf_min(cdf_min) );
  INV_X4 U1 ( .A(1'b1), .ZN(M2_WriteBus[36]) );
  INV_X4 U3 ( .A(1'b1), .ZN(M2_WriteBus[37]) );
  INV_X4 U5 ( .A(1'b1), .ZN(M2_WriteBus[38]) );
  INV_X4 U7 ( .A(1'b1), .ZN(M2_WriteBus[39]) );
  INV_X4 U9 ( .A(1'b1), .ZN(M2_WriteBus[40]) );
  INV_X4 U11 ( .A(1'b1), .ZN(M2_WriteBus[41]) );
  INV_X4 U13 ( .A(1'b1), .ZN(M2_WriteBus[42]) );
  INV_X4 U15 ( .A(1'b1), .ZN(M2_WriteBus[43]) );
  INV_X4 U17 ( .A(1'b1), .ZN(M2_WriteBus[44]) );
  INV_X4 U19 ( .A(1'b1), .ZN(M2_WriteBus[45]) );
  INV_X4 U21 ( .A(1'b1), .ZN(M2_WriteBus[46]) );
  INV_X4 U23 ( .A(1'b1), .ZN(M2_WriteBus[47]) );
  INV_X4 U25 ( .A(1'b1), .ZN(M2_WriteBus[48]) );
  INV_X4 U27 ( .A(1'b1), .ZN(M2_WriteBus[49]) );
  INV_X4 U29 ( .A(1'b1), .ZN(M2_WriteBus[50]) );
  INV_X4 U31 ( .A(1'b1), .ZN(M2_WriteBus[51]) );
  INV_X4 U33 ( .A(1'b1), .ZN(M2_WriteBus[52]) );
  INV_X4 U35 ( .A(1'b1), .ZN(M2_WriteBus[53]) );
  INV_X4 U37 ( .A(1'b1), .ZN(M2_WriteBus[54]) );
  INV_X4 U39 ( .A(1'b1), .ZN(M2_WriteBus[55]) );
  INV_X4 U41 ( .A(1'b1), .ZN(M2_WriteBus[56]) );
  INV_X4 U43 ( .A(1'b1), .ZN(M2_WriteBus[57]) );
  INV_X4 U45 ( .A(1'b1), .ZN(M2_WriteBus[58]) );
  INV_X4 U47 ( .A(1'b1), .ZN(M2_WriteBus[59]) );
  INV_X4 U49 ( .A(1'b1), .ZN(M2_WriteBus[60]) );
  INV_X4 U51 ( .A(1'b1), .ZN(M2_WriteBus[61]) );
  INV_X4 U53 ( .A(1'b1), .ZN(M2_WriteBus[62]) );
  INV_X4 U55 ( .A(1'b1), .ZN(M2_WriteBus[63]) );
  INV_X4 U57 ( .A(1'b1), .ZN(M2_WriteBus[64]) );
  INV_X4 U59 ( .A(1'b1), .ZN(M2_WriteBus[65]) );
  INV_X4 U61 ( .A(1'b1), .ZN(M2_WriteBus[66]) );
  INV_X4 U63 ( .A(1'b1), .ZN(M2_WriteBus[67]) );
  INV_X4 U65 ( .A(1'b1), .ZN(M2_WriteBus[68]) );
  INV_X4 U67 ( .A(1'b1), .ZN(M2_WriteBus[69]) );
  INV_X4 U69 ( .A(1'b1), .ZN(M2_WriteBus[70]) );
  INV_X4 U71 ( .A(1'b1), .ZN(M2_WriteBus[71]) );
  INV_X4 U73 ( .A(1'b1), .ZN(M2_WriteBus[72]) );
  INV_X4 U75 ( .A(1'b1), .ZN(M2_WriteBus[73]) );
  INV_X4 U77 ( .A(1'b1), .ZN(M2_WriteBus[74]) );
  INV_X4 U79 ( .A(1'b1), .ZN(M2_WriteBus[75]) );
  INV_X4 U81 ( .A(1'b1), .ZN(M2_WriteBus[76]) );
  INV_X4 U83 ( .A(1'b1), .ZN(M2_WriteBus[77]) );
  INV_X4 U85 ( .A(1'b1), .ZN(M2_WriteBus[78]) );
  INV_X4 U87 ( .A(1'b1), .ZN(M2_WriteBus[79]) );
  INV_X4 U89 ( .A(1'b1), .ZN(M2_WriteBus[80]) );
  INV_X4 U91 ( .A(1'b1), .ZN(M2_WriteBus[81]) );
  INV_X4 U93 ( .A(1'b1), .ZN(M2_WriteBus[82]) );
  INV_X4 U95 ( .A(1'b1), .ZN(M2_WriteBus[83]) );
  INV_X4 U97 ( .A(1'b1), .ZN(M2_WriteBus[84]) );
  INV_X4 U99 ( .A(1'b1), .ZN(M2_WriteBus[85]) );
  INV_X4 U101 ( .A(1'b1), .ZN(M2_WriteBus[86]) );
  INV_X4 U103 ( .A(1'b1), .ZN(M2_WriteBus[87]) );
  INV_X4 U105 ( .A(1'b1), .ZN(M2_WriteBus[88]) );
  INV_X4 U107 ( .A(1'b1), .ZN(M2_WriteBus[89]) );
  INV_X4 U109 ( .A(1'b1), .ZN(M2_WriteBus[90]) );
  INV_X4 U111 ( .A(1'b1), .ZN(M2_WriteBus[91]) );
  INV_X4 U113 ( .A(1'b1), .ZN(M2_WriteBus[92]) );
  INV_X4 U115 ( .A(1'b1), .ZN(M2_WriteBus[93]) );
  INV_X4 U117 ( .A(1'b1), .ZN(M2_WriteBus[94]) );
  INV_X4 U119 ( .A(1'b1), .ZN(M2_WriteBus[95]) );
  INV_X4 U121 ( .A(1'b1), .ZN(M2_WriteBus[96]) );
  INV_X4 U123 ( .A(1'b1), .ZN(M2_WriteBus[97]) );
  INV_X4 U125 ( .A(1'b1), .ZN(M2_WriteBus[98]) );
  INV_X4 U127 ( .A(1'b1), .ZN(M2_WriteBus[99]) );
  INV_X4 U129 ( .A(1'b1), .ZN(M2_WriteBus[100]) );
  INV_X4 U131 ( .A(1'b1), .ZN(M2_WriteBus[101]) );
  INV_X4 U133 ( .A(1'b1), .ZN(M2_WriteBus[102]) );
  INV_X4 U135 ( .A(1'b1), .ZN(M2_WriteBus[103]) );
  INV_X4 U137 ( .A(1'b1), .ZN(M2_WriteBus[104]) );
  INV_X4 U139 ( .A(1'b1), .ZN(M2_WriteBus[105]) );
  INV_X4 U141 ( .A(1'b1), .ZN(M2_WriteBus[106]) );
  INV_X4 U143 ( .A(1'b1), .ZN(M2_WriteBus[107]) );
  INV_X4 U145 ( .A(1'b1), .ZN(M2_WriteBus[108]) );
  INV_X4 U147 ( .A(1'b1), .ZN(M2_WriteBus[109]) );
  INV_X4 U149 ( .A(1'b1), .ZN(M2_WriteBus[110]) );
  INV_X4 U151 ( .A(1'b1), .ZN(M2_WriteBus[111]) );
  INV_X4 U153 ( .A(1'b1), .ZN(M2_WriteBus[112]) );
  INV_X4 U155 ( .A(1'b1), .ZN(M2_WriteBus[113]) );
  INV_X4 U157 ( .A(1'b1), .ZN(M2_WriteBus[114]) );
  INV_X4 U159 ( .A(1'b1), .ZN(M2_WriteBus[115]) );
  INV_X4 U161 ( .A(1'b1), .ZN(M2_WriteBus[116]) );
  INV_X4 U163 ( .A(1'b1), .ZN(M2_WriteBus[117]) );
  INV_X4 U165 ( .A(1'b1), .ZN(M2_WriteBus[118]) );
  INV_X4 U167 ( .A(1'b1), .ZN(M2_WriteBus[119]) );
  INV_X4 U169 ( .A(1'b1), .ZN(M2_WriteBus[120]) );
  INV_X4 U171 ( .A(1'b1), .ZN(M2_WriteBus[121]) );
  INV_X4 U173 ( .A(1'b1), .ZN(M2_WriteBus[122]) );
  INV_X4 U175 ( .A(1'b1), .ZN(M2_WriteBus[123]) );
  INV_X4 U177 ( .A(1'b1), .ZN(M2_WriteBus[124]) );
  INV_X4 U179 ( .A(1'b1), .ZN(M2_WriteBus[125]) );
  INV_X4 U181 ( .A(1'b1), .ZN(M2_WriteBus[126]) );
  INV_X4 U183 ( .A(1'b1), .ZN(M2_WriteBus[127]) );
  INV_X4 U185 ( .A(1'b1), .ZN(M2_ReadAddress2[8]) );
  INV_X4 U187 ( .A(1'b1), .ZN(M2_ReadAddress2[9]) );
  INV_X4 U189 ( .A(1'b1), .ZN(M2_ReadAddress2[10]) );
  INV_X4 U191 ( .A(1'b1), .ZN(M2_ReadAddress2[11]) );
  INV_X4 U193 ( .A(1'b1), .ZN(M2_ReadAddress2[12]) );
  INV_X4 U195 ( .A(1'b1), .ZN(M2_ReadAddress2[13]) );
  INV_X4 U197 ( .A(1'b1), .ZN(M2_ReadAddress2[14]) );
  INV_X4 U199 ( .A(n201), .ZN(n200) );
  INV_X4 U200 ( .A(reset_n), .ZN(n201) );
endmodule


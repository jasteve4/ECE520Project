
module Output_Fetch_MEM ( clock, reset_n, start, ReadBus, ReadAddress, DataOut, 
        StartOut, output_base_offset, done );
  input [127:0] ReadBus;
  output [15:0] ReadAddress;
  output [15:0] DataOut;
  input clock, reset_n, start, output_base_offset;
  output StartOut, done;
  wire   n415, n417, n418, n419, n420, n421, n422, n423, n424, \U3/U1/DATA1_0 ,
         \U3/U1/DATA1_1 , \U3/U1/DATA1_2 , \U3/U1/DATA1_3 , \U3/U1/DATA1_4 ,
         \U3/U1/DATA1_5 , \U3/U1/DATA1_6 , \U3/U1/DATA1_7 , \U3/U1/DATA1_8 ,
         \U3/U1/DATA1_9 , \U3/U1/DATA1_10 , \U3/U1/DATA1_11 , \U3/U1/DATA1_12 ,
         \U3/U1/DATA1_13 , \U3/U1/DATA1_14 , \U3/U1/DATA1_15 ,
         \U3/U1/DATA1_16 , \U3/U1/DATA1_17 , \U3/U1/DATA1_18 ,
         \U3/U1/DATA1_19 , \U3/U1/DATA1_20 , \U3/U1/DATA1_21 ,
         \U3/U1/DATA1_22 , \U3/U1/DATA1_23 , \U3/U1/DATA1_24 ,
         \U3/U1/DATA1_25 , \U3/U1/DATA1_26 , \U3/U1/DATA1_27 ,
         \U3/U1/DATA1_28 , \U3/U1/DATA1_29 , \U3/U1/DATA1_30 ,
         \U3/U1/DATA1_31 , \U3/U1/DATA1_32 , \U3/U1/DATA1_33 ,
         \U3/U1/DATA1_34 , \U3/U1/DATA1_35 , \U3/U1/DATA1_36 ,
         \U3/U1/DATA1_37 , \U3/U1/DATA1_38 , \U3/U1/DATA1_39 ,
         \U3/U1/DATA1_40 , \U3/U1/DATA1_41 , \U3/U1/DATA1_42 ,
         \U3/U1/DATA1_43 , \U3/U1/DATA1_44 , \U3/U1/DATA1_45 ,
         \U3/U1/DATA1_46 , \U3/U1/DATA1_47 , \U3/U1/DATA1_48 ,
         \U3/U1/DATA1_49 , \U3/U1/DATA1_50 , \U3/U1/DATA1_51 ,
         \U3/U1/DATA1_52 , \U3/U1/DATA1_53 , \U3/U1/DATA1_54 ,
         \U3/U1/DATA1_55 , \U3/U1/DATA1_56 , \U3/U1/DATA1_57 ,
         \U3/U1/DATA1_58 , \U3/U1/DATA1_59 , \U3/U1/DATA1_60 ,
         \U3/U1/DATA1_61 , \U3/U1/DATA1_62 , \U3/U1/DATA1_63 ,
         \U3/U1/DATA1_64 , \U3/U1/DATA1_65 , \U3/U1/DATA1_66 ,
         \U3/U1/DATA1_67 , \U3/U1/DATA1_68 , \U3/U1/DATA1_69 ,
         \U3/U1/DATA1_70 , \U3/U1/DATA1_71 , \U3/U1/DATA1_72 ,
         \U3/U1/DATA1_73 , \U3/U1/DATA1_74 , \U3/U1/DATA1_75 ,
         \U3/U1/DATA1_76 , \U3/U1/DATA1_77 , \U3/U1/DATA1_78 ,
         \U3/U1/DATA1_79 , \U3/U1/DATA1_80 , \U3/U1/DATA1_81 ,
         \U3/U1/DATA1_82 , \U3/U1/DATA1_83 , \U3/U1/DATA1_84 ,
         \U3/U1/DATA1_85 , \U3/U1/DATA1_86 , \U3/U1/DATA1_87 ,
         \U3/U1/DATA1_88 , \U3/U1/DATA1_89 , \U3/U1/DATA1_90 ,
         \U3/U1/DATA1_91 , \U3/U1/DATA1_92 , \U3/U1/DATA1_93 ,
         \U3/U1/DATA1_94 , \U3/U1/DATA1_95 , \U3/U1/DATA1_96 ,
         \U3/U1/DATA1_97 , \U3/U1/DATA1_98 , \U3/U1/DATA1_99 ,
         \U3/U1/DATA1_100 , \U3/U1/DATA1_101 , \U3/U1/DATA1_102 ,
         \U3/U1/DATA1_103 , \U3/U1/DATA1_104 , \U3/U1/DATA1_105 ,
         \U3/U1/DATA1_106 , \U3/U1/DATA1_107 , \U3/U1/DATA1_108 ,
         \U3/U1/DATA1_109 , \U3/U1/DATA1_110 , \U3/U1/DATA1_111 ,
         \U3/U1/DATA1_112 , \U3/U1/DATA1_113 , \U3/U1/DATA1_114 ,
         \U3/U1/DATA1_115 , \U3/U1/DATA1_116 , \U3/U1/DATA1_117 ,
         \U3/U1/DATA1_118 , \U3/U1/DATA1_119 , \U3/U2/DATA2_15 , \U3/U3/Z_0 ,
         \U3/U4/Z_0 , \U3/U5/Z_0 , \U3/U5/Z_1 , \U3/U5/Z_2 , \U3/U5/Z_3 ,
         \U6/DATA1_0 , \U6/DATA1_1 , \U6/DATA1_2 , \U6/DATA1_3 , \U5/Z_0 ,
         \U5/Z_1 , \U5/Z_2 , \U5/Z_3 , \U5/Z_4 , \U5/Z_5 , \U5/Z_6 , \U5/Z_7 ,
         \U5/DATA16_0 , \U5/DATA16_1 , \U5/DATA16_2 , \U5/DATA16_3 ,
         \U5/DATA16_4 , \U5/DATA16_5 , \U5/DATA16_6 , \U5/DATA16_7 ,
         \U5/DATA15_0 , \U5/DATA15_1 , \U5/DATA15_2 , \U5/DATA15_3 ,
         \U5/DATA15_4 , \U5/DATA15_5 , \U5/DATA15_6 , \U5/DATA15_7 ,
         \U5/DATA14_0 , \U5/DATA14_1 , \U5/DATA14_2 , \U5/DATA14_3 ,
         \U5/DATA14_4 , \U5/DATA14_5 , \U5/DATA14_6 , \U5/DATA14_7 ,
         \U5/DATA13_0 , \U5/DATA13_1 , \U5/DATA13_2 , \U5/DATA13_3 ,
         \U5/DATA13_4 , \U5/DATA13_5 , \U5/DATA13_6 , \U5/DATA13_7 ,
         \U5/DATA12_0 , \U5/DATA12_1 , \U5/DATA12_2 , \U5/DATA12_3 ,
         \U5/DATA12_4 , \U5/DATA12_5 , \U5/DATA12_6 , \U5/DATA12_7 ,
         \U5/DATA11_0 , \U5/DATA11_1 , \U5/DATA11_2 , \U5/DATA11_3 ,
         \U5/DATA11_4 , \U5/DATA11_5 , \U5/DATA11_6 , \U5/DATA11_7 ,
         \U5/DATA10_0 , \U5/DATA10_1 , \U5/DATA10_2 , \U5/DATA10_3 ,
         \U5/DATA10_4 , \U5/DATA10_5 , \U5/DATA10_6 , \U5/DATA10_7 ,
         \U5/DATA9_0 , \U5/DATA9_1 , \U5/DATA9_2 , \U5/DATA9_3 , \U5/DATA9_4 ,
         \U5/DATA9_5 , \U5/DATA9_6 , \U5/DATA9_7 , \U5/DATA8_0 , \U5/DATA8_1 ,
         \U5/DATA8_2 , \U5/DATA8_3 , \U5/DATA8_4 , \U5/DATA8_5 , \U5/DATA8_6 ,
         \U5/DATA8_7 , \U5/DATA7_0 , \U5/DATA7_1 , \U5/DATA7_2 , \U5/DATA7_3 ,
         \U5/DATA7_4 , \U5/DATA7_5 , \U5/DATA7_6 , \U5/DATA7_7 , \U5/DATA6_0 ,
         \U5/DATA6_1 , \U5/DATA6_2 , \U5/DATA6_3 , \U5/DATA6_4 , \U5/DATA6_5 ,
         \U5/DATA6_6 , \U5/DATA6_7 , \U5/DATA5_0 , \U5/DATA5_1 , \U5/DATA5_2 ,
         \U5/DATA5_3 , \U5/DATA5_4 , \U5/DATA5_5 , \U5/DATA5_6 , \U5/DATA5_7 ,
         \U5/DATA4_0 , \U5/DATA4_1 , \U5/DATA4_2 , \U5/DATA4_3 , \U5/DATA4_4 ,
         \U5/DATA4_5 , \U5/DATA4_6 , \U5/DATA4_7 , \U5/DATA3_0 , \U5/DATA3_1 ,
         \U5/DATA3_2 , \U5/DATA3_3 , \U5/DATA3_4 , \U5/DATA3_5 , \U5/DATA3_6 ,
         \U5/DATA3_7 , \U5/DATA2_0 , \U5/DATA2_1 , \U5/DATA2_2 , \U5/DATA2_3 ,
         \U5/DATA2_4 , \U5/DATA2_5 , \U5/DATA2_6 , \U5/DATA2_7 , \U5/DATA1_0 ,
         \U5/DATA1_1 , \U5/DATA1_2 , \U5/DATA1_3 , \U5/DATA1_4 , \U5/DATA1_5 ,
         \U5/DATA1_6 , \U5/DATA1_7 , \U4/DATA1_0 , \U4/DATA1_1 , \U4/DATA1_2 ,
         \U4/DATA1_3 , \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 , \U4/DATA1_7 ,
         \U4/DATA1_8 , \U4/DATA1_9 , \U4/DATA1_10 , \U4/DATA1_11 ,
         \U4/DATA1_12 , \U4/DATA1_13 , \U4/DATA1_14 , \U4/DATA1_15 , n143,
         n145, n146, n147, n149, n155, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n280, n281,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727;
  assign \U3/U1/DATA1_0  = ReadBus[8];
  assign \U3/U1/DATA1_1  = ReadBus[9];
  assign \U3/U1/DATA1_2  = ReadBus[10];
  assign \U3/U1/DATA1_3  = ReadBus[11];
  assign \U3/U1/DATA1_4  = ReadBus[12];
  assign \U3/U1/DATA1_5  = ReadBus[13];
  assign \U3/U1/DATA1_6  = ReadBus[14];
  assign \U3/U1/DATA1_7  = ReadBus[15];
  assign \U3/U1/DATA1_8  = ReadBus[16];
  assign \U3/U1/DATA1_9  = ReadBus[17];
  assign \U3/U1/DATA1_10  = ReadBus[18];
  assign \U3/U1/DATA1_11  = ReadBus[19];
  assign \U3/U1/DATA1_12  = ReadBus[20];
  assign \U3/U1/DATA1_13  = ReadBus[21];
  assign \U3/U1/DATA1_14  = ReadBus[22];
  assign \U3/U1/DATA1_15  = ReadBus[23];
  assign \U3/U1/DATA1_16  = ReadBus[24];
  assign \U3/U1/DATA1_17  = ReadBus[25];
  assign \U3/U1/DATA1_18  = ReadBus[26];
  assign \U3/U1/DATA1_19  = ReadBus[27];
  assign \U3/U1/DATA1_20  = ReadBus[28];
  assign \U3/U1/DATA1_21  = ReadBus[29];
  assign \U3/U1/DATA1_22  = ReadBus[30];
  assign \U3/U1/DATA1_23  = ReadBus[31];
  assign \U3/U1/DATA1_24  = ReadBus[32];
  assign \U3/U1/DATA1_25  = ReadBus[33];
  assign \U3/U1/DATA1_26  = ReadBus[34];
  assign \U3/U1/DATA1_27  = ReadBus[35];
  assign \U3/U1/DATA1_28  = ReadBus[36];
  assign \U3/U1/DATA1_29  = ReadBus[37];
  assign \U3/U1/DATA1_30  = ReadBus[38];
  assign \U3/U1/DATA1_31  = ReadBus[39];
  assign \U3/U1/DATA1_32  = ReadBus[40];
  assign \U3/U1/DATA1_33  = ReadBus[41];
  assign \U3/U1/DATA1_34  = ReadBus[42];
  assign \U3/U1/DATA1_35  = ReadBus[43];
  assign \U3/U1/DATA1_36  = ReadBus[44];
  assign \U3/U1/DATA1_37  = ReadBus[45];
  assign \U3/U1/DATA1_38  = ReadBus[46];
  assign \U3/U1/DATA1_39  = ReadBus[47];
  assign \U3/U1/DATA1_40  = ReadBus[48];
  assign \U3/U1/DATA1_41  = ReadBus[49];
  assign \U3/U1/DATA1_42  = ReadBus[50];
  assign \U3/U1/DATA1_43  = ReadBus[51];
  assign \U3/U1/DATA1_44  = ReadBus[52];
  assign \U3/U1/DATA1_45  = ReadBus[53];
  assign \U3/U1/DATA1_46  = ReadBus[54];
  assign \U3/U1/DATA1_47  = ReadBus[55];
  assign \U3/U1/DATA1_48  = ReadBus[56];
  assign \U3/U1/DATA1_49  = ReadBus[57];
  assign \U3/U1/DATA1_50  = ReadBus[58];
  assign \U3/U1/DATA1_51  = ReadBus[59];
  assign \U3/U1/DATA1_52  = ReadBus[60];
  assign \U3/U1/DATA1_53  = ReadBus[61];
  assign \U3/U1/DATA1_54  = ReadBus[62];
  assign \U3/U1/DATA1_55  = ReadBus[63];
  assign \U3/U1/DATA1_56  = ReadBus[64];
  assign \U3/U1/DATA1_57  = ReadBus[65];
  assign \U3/U1/DATA1_58  = ReadBus[66];
  assign \U3/U1/DATA1_59  = ReadBus[67];
  assign \U3/U1/DATA1_60  = ReadBus[68];
  assign \U3/U1/DATA1_61  = ReadBus[69];
  assign \U3/U1/DATA1_62  = ReadBus[70];
  assign \U3/U1/DATA1_63  = ReadBus[71];
  assign \U3/U1/DATA1_64  = ReadBus[72];
  assign \U3/U1/DATA1_65  = ReadBus[73];
  assign \U3/U1/DATA1_66  = ReadBus[74];
  assign \U3/U1/DATA1_67  = ReadBus[75];
  assign \U3/U1/DATA1_68  = ReadBus[76];
  assign \U3/U1/DATA1_69  = ReadBus[77];
  assign \U3/U1/DATA1_70  = ReadBus[78];
  assign \U3/U1/DATA1_71  = ReadBus[79];
  assign \U3/U1/DATA1_72  = ReadBus[80];
  assign \U3/U1/DATA1_73  = ReadBus[81];
  assign \U3/U1/DATA1_74  = ReadBus[82];
  assign \U3/U1/DATA1_75  = ReadBus[83];
  assign \U3/U1/DATA1_76  = ReadBus[84];
  assign \U3/U1/DATA1_77  = ReadBus[85];
  assign \U3/U1/DATA1_78  = ReadBus[86];
  assign \U3/U1/DATA1_79  = ReadBus[87];
  assign \U3/U1/DATA1_80  = ReadBus[88];
  assign \U3/U1/DATA1_81  = ReadBus[89];
  assign \U3/U1/DATA1_82  = ReadBus[90];
  assign \U3/U1/DATA1_83  = ReadBus[91];
  assign \U3/U1/DATA1_84  = ReadBus[92];
  assign \U3/U1/DATA1_85  = ReadBus[93];
  assign \U3/U1/DATA1_86  = ReadBus[94];
  assign \U3/U1/DATA1_87  = ReadBus[95];
  assign \U3/U1/DATA1_88  = ReadBus[96];
  assign \U3/U1/DATA1_89  = ReadBus[97];
  assign \U3/U1/DATA1_90  = ReadBus[98];
  assign \U3/U1/DATA1_91  = ReadBus[99];
  assign \U3/U1/DATA1_92  = ReadBus[100];
  assign \U3/U1/DATA1_93  = ReadBus[101];
  assign \U3/U1/DATA1_94  = ReadBus[102];
  assign \U3/U1/DATA1_95  = ReadBus[103];
  assign \U3/U1/DATA1_96  = ReadBus[104];
  assign \U3/U1/DATA1_97  = ReadBus[105];
  assign \U3/U1/DATA1_98  = ReadBus[106];
  assign \U3/U1/DATA1_99  = ReadBus[107];
  assign \U3/U1/DATA1_100  = ReadBus[108];
  assign \U3/U1/DATA1_101  = ReadBus[109];
  assign \U3/U1/DATA1_102  = ReadBus[110];
  assign \U3/U1/DATA1_103  = ReadBus[111];
  assign \U3/U1/DATA1_104  = ReadBus[112];
  assign \U3/U1/DATA1_105  = ReadBus[113];
  assign \U3/U1/DATA1_106  = ReadBus[114];
  assign \U3/U1/DATA1_107  = ReadBus[115];
  assign \U3/U1/DATA1_108  = ReadBus[116];
  assign \U3/U1/DATA1_109  = ReadBus[117];
  assign \U3/U1/DATA1_110  = ReadBus[118];
  assign \U3/U1/DATA1_111  = ReadBus[119];
  assign \U3/U1/DATA1_112  = ReadBus[120];
  assign \U3/U1/DATA1_113  = ReadBus[121];
  assign \U3/U1/DATA1_114  = ReadBus[122];
  assign \U3/U1/DATA1_115  = ReadBus[123];
  assign \U3/U1/DATA1_116  = ReadBus[124];
  assign \U3/U1/DATA1_117  = ReadBus[125];
  assign \U3/U1/DATA1_118  = ReadBus[126];
  assign \U3/U1/DATA1_119  = ReadBus[127];
  assign \U3/U2/DATA2_15  = output_base_offset;
  assign DataOut[0] = \U5/Z_0 ;
  assign DataOut[1] = \U5/Z_1 ;
  assign DataOut[2] = \U5/Z_2 ;
  assign DataOut[3] = \U5/Z_3 ;
  assign DataOut[4] = \U5/Z_4 ;
  assign DataOut[5] = \U5/Z_5 ;
  assign DataOut[6] = \U5/Z_6 ;
  assign DataOut[7] = \U5/Z_7 ;
  assign ReadAddress[0] = \U4/DATA1_0 ;
  assign ReadAddress[1] = \U4/DATA1_1 ;
  assign ReadAddress[2] = \U4/DATA1_2 ;
  assign ReadAddress[3] = \U4/DATA1_3 ;
  assign ReadAddress[4] = \U4/DATA1_4 ;
  assign ReadAddress[5] = \U4/DATA1_5 ;
  assign ReadAddress[6] = \U4/DATA1_6 ;
  assign ReadAddress[7] = \U4/DATA1_7 ;
  assign ReadAddress[8] = \U4/DATA1_8 ;
  assign ReadAddress[9] = \U4/DATA1_9 ;
  assign ReadAddress[10] = \U4/DATA1_10 ;
  assign ReadAddress[11] = \U4/DATA1_11 ;
  assign ReadAddress[12] = \U4/DATA1_12 ;
  assign ReadAddress[13] = \U4/DATA1_13 ;
  assign ReadAddress[14] = \U4/DATA1_14 ;
  assign ReadAddress[15] = \U4/DATA1_15 ;

  DFF_X1 \data_in_reg[7]  ( .D(ReadBus[7]), .CK(clock), .Q(\U5/DATA16_7 ) );
  DFF_X1 \data_in_reg[6]  ( .D(ReadBus[6]), .CK(clock), .Q(\U5/DATA16_6 ) );
  DFF_X1 \data_in_reg[5]  ( .D(ReadBus[5]), .CK(clock), .Q(\U5/DATA16_5 ) );
  DFF_X1 \data_in_reg[4]  ( .D(ReadBus[4]), .CK(clock), .Q(\U5/DATA16_4 ) );
  DFF_X1 \data_in_reg[3]  ( .D(ReadBus[3]), .CK(clock), .Q(\U5/DATA16_3 ) );
  DFF_X1 \data_in_reg[2]  ( .D(ReadBus[2]), .CK(clock), .Q(\U5/DATA16_2 ) );
  DFF_X1 \data_in_reg[1]  ( .D(ReadBus[1]), .CK(clock), .Q(\U5/DATA16_1 ) );
  DFF_X1 \data_in_reg[0]  ( .D(ReadBus[0]), .CK(clock), .Q(\U5/DATA16_0 ) );
  SDFFR_X2 \data_in_reg[107]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_99 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA13_3 ) );
  SDFFR_X2 \data_in_reg[106]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_98 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA13_2 ) );
  SDFFR_X2 \data_in_reg[105]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_97 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA13_1 ) );
  SDFFR_X2 \data_in_reg[104]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_96 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA13_0 ) );
  SDFFR_X2 \data_in_reg[103]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_95 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA12_7 ) );
  SDFFR_X2 \data_in_reg[102]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_94 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA12_6 ) );
  SDFFR_X2 \data_in_reg[101]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_93 ), 
        .CK(clock), .RN(n623), .Q(\U5/DATA12_5 ) );
  SDFFR_X2 \data_in_reg[100]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_92 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA12_4 ) );
  SDFFR_X2 \data_in_reg[99]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_91 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA12_3 ) );
  SDFFR_X2 \data_in_reg[98]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_90 ), 
        .CK(clock), .RN(n623), .Q(\U5/DATA12_2 ) );
  SDFFR_X2 \data_in_reg[17]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_9 ), .CK(
        clock), .RN(n624), .Q(\U5/DATA2_1 ) );
  SDFFR_X2 \data_in_reg[97]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_89 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA12_1 ) );
  SDFFR_X2 \data_in_reg[96]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_88 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA12_0 ) );
  SDFFR_X2 \data_in_reg[95]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_87 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA11_7 ) );
  SDFFR_X2 \data_in_reg[94]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_86 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA11_6 ) );
  SDFFR_X2 \data_in_reg[93]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_85 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA11_5 ) );
  SDFFR_X2 \data_in_reg[92]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_84 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA11_4 ) );
  SDFFR_X2 \data_in_reg[91]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_83 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA11_3 ) );
  SDFFR_X2 \data_in_reg[90]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_82 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA11_2 ) );
  SDFFR_X2 \data_in_reg[89]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_81 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA11_1 ) );
  SDFFR_X2 \data_in_reg[88]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_80 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA11_0 ) );
  SDFFR_X2 \data_in_reg[16]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_8 ), .CK(
        clock), .RN(n624), .Q(\U5/DATA2_0 ) );
  SDFFR_X2 \data_in_reg[87]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_79 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA10_7 ) );
  SDFFR_X2 \data_in_reg[86]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_78 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA10_6 ) );
  SDFFR_X2 \data_in_reg[85]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_77 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA10_5 ) );
  SDFFR_X2 \data_in_reg[84]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_76 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA10_4 ) );
  SDFFR_X2 \data_in_reg[83]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_75 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA10_3 ) );
  SDFFR_X2 \data_in_reg[82]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_74 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA10_2 ) );
  SDFFR_X2 \data_in_reg[81]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_73 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA10_1 ) );
  SDFFR_X2 \data_in_reg[80]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_72 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA10_0 ) );
  SDFFR_X2 \data_in_reg[79]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_71 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA9_7 ) );
  SDFFR_X2 \data_in_reg[78]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_70 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA9_6 ) );
  SDFFR_X2 \data_in_reg[15]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_7 ), .CK(
        clock), .RN(n624), .Q(\U5/DATA1_7 ) );
  SDFFR_X2 \data_in_reg[77]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_69 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA9_5 ) );
  SDFFR_X2 \data_in_reg[76]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_68 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA9_4 ) );
  SDFFR_X2 \data_in_reg[75]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_67 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA9_3 ) );
  SDFFR_X2 \data_in_reg[74]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_66 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA9_2 ) );
  SDFFR_X2 \data_in_reg[73]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_65 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA9_1 ) );
  SDFFR_X2 \data_in_reg[72]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_64 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA9_0 ) );
  SDFFR_X2 \data_in_reg[71]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_63 ), 
        .CK(clock), .RN(n624), .Q(\U5/DATA8_7 ) );
  SDFFR_X2 \data_in_reg[70]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_62 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA8_6 ) );
  SDFFR_X2 \data_in_reg[69]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_61 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA8_5 ) );
  SDFFR_X2 \data_in_reg[68]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_60 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA8_4 ) );
  SDFFR_X2 \data_in_reg[14]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_6 ), .CK(
        clock), .RN(n625), .Q(\U5/DATA1_6 ) );
  SDFFR_X2 \data_in_reg[67]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_59 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA8_3 ) );
  SDFFR_X2 \data_in_reg[66]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_58 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA8_2 ) );
  SDFFR_X2 \data_in_reg[65]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_57 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA8_1 ) );
  SDFFR_X2 \data_in_reg[64]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_56 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA8_0 ) );
  SDFFR_X2 \data_in_reg[63]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_55 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA7_7 ) );
  SDFFR_X2 \data_in_reg[62]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_54 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA7_6 ) );
  SDFFR_X2 \data_in_reg[61]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_53 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA7_5 ) );
  SDFFR_X2 \data_in_reg[60]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_52 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA7_4 ) );
  SDFFR_X2 \data_in_reg[59]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_51 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA7_3 ) );
  SDFFR_X2 \data_in_reg[58]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_50 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA7_2 ) );
  SDFFR_X2 \data_in_reg[13]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_5 ), .CK(
        clock), .RN(n625), .Q(\U5/DATA1_5 ) );
  SDFFR_X2 \data_in_reg[57]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_49 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA7_1 ) );
  SDFFR_X2 \data_in_reg[56]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_48 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA7_0 ) );
  SDFFR_X2 \data_in_reg[55]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_47 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA6_7 ) );
  SDFFR_X2 \data_in_reg[54]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_46 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA6_6 ) );
  SDFFR_X2 \data_in_reg[53]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_45 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA6_5 ) );
  SDFFR_X2 \data_in_reg[52]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_44 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA6_4 ) );
  SDFFR_X2 \data_in_reg[51]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_43 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA6_3 ) );
  SDFFR_X2 \data_in_reg[50]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_42 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA6_2 ) );
  SDFFR_X2 \data_in_reg[49]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_41 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA6_1 ) );
  SDFFR_X2 \data_in_reg[48]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_40 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA6_0 ) );
  SDFFR_X2 \data_in_reg[12]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_4 ), .CK(
        clock), .RN(n625), .Q(\U5/DATA1_4 ) );
  SDFFR_X2 \data_in_reg[47]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_39 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA5_7 ) );
  SDFFR_X2 \data_in_reg[46]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_38 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA5_6 ) );
  SDFFR_X2 \data_in_reg[45]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_37 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA5_5 ) );
  SDFFR_X2 \data_in_reg[44]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_36 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA5_4 ) );
  SDFFR_X2 \data_in_reg[43]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_35 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA5_3 ) );
  SDFFR_X2 \data_in_reg[42]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_34 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA5_2 ) );
  SDFFR_X2 \data_in_reg[41]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_33 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA5_1 ) );
  SDFFR_X2 \data_in_reg[40]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_32 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA5_0 ) );
  SDFFR_X2 \data_in_reg[39]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_31 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA4_7 ) );
  SDFFR_X2 \data_in_reg[38]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_30 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA4_6 ) );
  SDFFR_X2 \data_in_reg[11]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_3 ), .CK(
        clock), .RN(n626), .Q(\U5/DATA1_3 ) );
  SDFFR_X2 \data_in_reg[37]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_29 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA4_5 ) );
  SDFFR_X2 \data_in_reg[36]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_28 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA4_4 ) );
  SDFFR_X2 \data_in_reg[35]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_27 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA4_3 ) );
  SDFFR_X2 \data_in_reg[34]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_26 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA4_2 ) );
  SDFFR_X2 \data_in_reg[33]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_25 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA4_1 ) );
  SDFFR_X2 \data_in_reg[32]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_24 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA4_0 ) );
  SDFFR_X2 \data_in_reg[31]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_23 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA3_7 ) );
  SDFFR_X2 \data_in_reg[30]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_22 ), 
        .CK(clock), .RN(n625), .Q(\U5/DATA3_6 ) );
  SDFFR_X2 \data_in_reg[29]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_21 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA3_5 ) );
  SDFFR_X2 \data_in_reg[28]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_20 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA3_4 ) );
  SDFFR_X2 \data_in_reg[10]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_2 ), .CK(
        clock), .RN(n626), .Q(\U5/DATA1_2 ) );
  SDFFR_X2 \data_in_reg[27]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_19 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA3_3 ) );
  SDFFR_X2 \data_in_reg[26]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_18 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA3_2 ) );
  SDFFR_X2 \data_in_reg[25]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_17 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA3_1 ) );
  SDFFR_X2 \data_in_reg[24]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_16 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA3_0 ) );
  SDFFR_X2 \data_in_reg[23]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_15 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA2_7 ) );
  SDFFR_X2 \data_in_reg[22]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_14 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA2_6 ) );
  SDFFR_X2 \data_in_reg[21]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_13 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA2_5 ) );
  SDFFR_X2 \data_in_reg[20]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_12 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA2_4 ) );
  SDFFR_X2 \data_in_reg[127]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_119 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA15_7 ) );
  SDFFR_X2 \data_in_reg[126]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_118 ), 
        .CK(clock), .RN(n626), .Q(\U5/DATA15_6 ) );
  SDFFR_X2 \data_in_reg[125]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_117 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA15_5 ) );
  SDFFR_X2 \data_in_reg[124]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_116 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA15_4 ) );
  SDFFR_X2 \data_in_reg[123]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_115 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA15_3 ) );
  SDFFR_X2 \data_in_reg[122]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_114 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA15_2 ) );
  SDFFR_X2 \data_in_reg[121]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_113 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA15_1 ) );
  SDFFR_X2 \data_in_reg[120]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_112 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA15_0 ) );
  SDFFR_X2 \data_in_reg[119]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_111 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA14_7 ) );
  SDFFR_X2 \data_in_reg[118]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_110 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA14_6 ) );
  SDFFR_X2 \data_in_reg[19]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_11 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA2_3 ) );
  SDFFR_X2 \data_in_reg[117]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_109 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA14_5 ) );
  SDFFR_X2 \data_in_reg[116]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_108 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA14_4 ) );
  SDFFR_X2 \data_in_reg[115]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_107 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA14_3 ) );
  SDFFR_X2 \data_in_reg[114]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_106 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA14_2 ) );
  SDFFR_X2 \data_in_reg[113]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_105 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA14_1 ) );
  SDFFR_X2 \data_in_reg[112]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_104 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA14_0 ) );
  SDFFR_X2 \data_in_reg[111]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_103 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA13_7 ) );
  SDFFR_X2 \data_in_reg[110]  ( .D(1'b0), .SI(n620), .SE(\U3/U1/DATA1_102 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA13_6 ) );
  SDFFR_X2 \data_in_reg[109]  ( .D(1'b0), .SI(start), .SE(\U3/U1/DATA1_101 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA13_5 ) );
  SDFFR_X2 \data_in_reg[108]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_100 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA13_4 ) );
  SDFFR_X2 \data_in_reg[18]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_10 ), 
        .CK(clock), .RN(n627), .Q(\U5/DATA2_2 ) );
  SDFFR_X2 \data_in_reg[9]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_1 ), .CK(
        clock), .RN(n627), .Q(\U5/DATA1_1 ) );
  SDFFR_X2 \data_in_reg[8]  ( .D(1'b0), .SI(n619), .SE(\U3/U1/DATA1_0 ), .CK(
        clock), .RN(n623), .Q(\U5/DATA1_0 ) );
  NAND4_X2 U143 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(n174) );
  NAND4_X2 U148 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(n173) );
  NAND4_X2 U153 ( .A1(n201), .A2(n202), .A3(n203), .A4(n204), .ZN(n200) );
  NAND4_X2 U158 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(n199) );
  NAND4_X2 U163 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(n210) );
  NAND4_X2 U168 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(n209) );
  NAND4_X2 U173 ( .A1(n221), .A2(n222), .A3(n223), .A4(n224), .ZN(n220) );
  NAND4_X2 U178 ( .A1(n225), .A2(n226), .A3(n227), .A4(n228), .ZN(n219) );
  NAND4_X2 U183 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(n230) );
  NAND4_X2 U188 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(n229) );
  NAND4_X2 U193 ( .A1(n241), .A2(n242), .A3(n243), .A4(n244), .ZN(n240) );
  NAND4_X2 U198 ( .A1(n245), .A2(n246), .A3(n247), .A4(n248), .ZN(n239) );
  NAND4_X2 U203 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(n250) );
  NAND4_X2 U208 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(n249) );
  NAND4_X2 U213 ( .A1(n261), .A2(n262), .A3(n263), .A4(n264), .ZN(n260) );
  NOR3_X2 U215 ( .A1(n143), .A2(\U6/DATA1_2 ), .A3(n265), .ZN(n180) );
  NOR4_X2 U216 ( .A1(n143), .A2(\U6/DATA1_0 ), .A3(\U6/DATA1_1 ), .A4(
        \U6/DATA1_2 ), .ZN(n179) );
  AND3_X2 U218 ( .A1(\U6/DATA1_3 ), .A2(\U6/DATA1_0 ), .A3(n618), .ZN(n182) );
  AND3_X2 U219 ( .A1(\U6/DATA1_3 ), .A2(n146), .A3(n618), .ZN(n181) );
  NOR3_X2 U221 ( .A1(n143), .A2(n707), .A3(n265), .ZN(n184) );
  AND3_X2 U222 ( .A1(\U6/DATA1_3 ), .A2(n145), .A3(n267), .ZN(n183) );
  AND3_X2 U224 ( .A1(\U6/DATA1_3 ), .A2(\U6/DATA1_1 ), .A3(n267), .ZN(n185) );
  NAND4_X2 U225 ( .A1(n268), .A2(n269), .A3(n270), .A4(n271), .ZN(n259) );
  NOR3_X2 U227 ( .A1(\U6/DATA1_2 ), .A2(\U6/DATA1_3 ), .A3(n265), .ZN(n192) );
  NOR4_X2 U228 ( .A1(\U6/DATA1_0 ), .A2(\U6/DATA1_1 ), .A3(\U6/DATA1_2 ), .A4(
        \U6/DATA1_3 ), .ZN(n191) );
  AND3_X2 U230 ( .A1(\U6/DATA1_0 ), .A2(n143), .A3(n618), .ZN(n194) );
  AND3_X2 U231 ( .A1(n146), .A2(n143), .A3(n618), .ZN(n193) );
  NOR3_X2 U233 ( .A1(n707), .A2(\U6/DATA1_3 ), .A3(n265), .ZN(n196) );
  AND3_X2 U234 ( .A1(n145), .A2(n143), .A3(n267), .ZN(n195) );
  AND3_X2 U236 ( .A1(\U6/DATA1_1 ), .A2(n143), .A3(n267), .ZN(n197) );
  NOR2_X2 U237 ( .A1(n707), .A2(\U6/DATA1_0 ), .ZN(n267) );
  NOR4_X2 U240 ( .A1(n707), .A2(n145), .A3(n146), .A4(\U6/DATA1_3 ), .ZN(n198)
         );
  OAI22_X2 U245 ( .A1(n265), .A2(n172), .B1(n275), .B2(n145), .ZN(\U3/U5/Z_1 )
         );
  NAND2_X2 U247 ( .A1(\U6/DATA1_0 ), .A2(n145), .ZN(n265) );
  NOR2_X2 U249 ( .A1(n171), .A2(n155), .ZN(\U3/U4/Z_0 ) );
  DFFR_X2 \short_count_reg[3]  ( .D(\U3/U5/Z_3 ), .CK(clock), .RN(n622), .Q(
        \U6/DATA1_3 ), .QN(n143) );
  DFFR_X2 \ReadAddress_reg[15]  ( .D(n280), .CK(clock), .RN(n622), .Q(
        \U4/DATA1_15 ), .QN(n147) );
  DFFR_X2 \ReadAddress_reg[0]  ( .D(n281), .CK(clock), .RN(reset_n), .Q(
        \U4/DATA1_0 ), .QN(n149) );
  DFF_X2 base_offset_reg ( .D(\U3/U2/DATA2_15 ), .CK(clock), .Q(DataOut[15])
         );
  DFFR_X2 \short_count_reg[0]  ( .D(\U3/U5/Z_0 ), .CK(clock), .RN(n623), .Q(
        \U6/DATA1_0 ), .QN(n146) );
  DFFR_X2 \short_count_reg[1]  ( .D(\U3/U5/Z_1 ), .CK(clock), .RN(n623), .Q(
        \U6/DATA1_1 ), .QN(n145) );
  DFFR_X2 \short_count_reg[2]  ( .D(\U3/U5/Z_2 ), .CK(clock), .RN(n623), .Q(
        \U6/DATA1_2 ), .QN(n707) );
  DFFR_X2 done_reg ( .D(n415), .CK(clock), .RN(n622), .Q(done) );
  DFFR_X2 done8_reg ( .D(n417), .CK(clock), .RN(n622), .Q(n415) );
  DFFR_X2 done7_reg ( .D(n418), .CK(clock), .RN(n622), .Q(n417) );
  DFFR_X2 done6_reg ( .D(n419), .CK(clock), .RN(n622), .Q(n418) );
  DFFR_X2 done5_reg ( .D(n420), .CK(clock), .RN(n622), .Q(n419) );
  DFFR_X2 done4_reg ( .D(n421), .CK(clock), .RN(n622), .Q(n420) );
  DFFR_X2 done3_reg ( .D(n422), .CK(clock), .RN(n622), .Q(n421) );
  DFFR_X2 done2_reg ( .D(n423), .CK(clock), .RN(n622), .Q(n422) );
  DFFR_X2 done1_reg ( .D(n424), .CK(clock), .RN(n622), .Q(n423) );
  DFFR_X2 StartOut_reg ( .D(\U3/U3/Z_0 ), .CK(clock), .RN(reset_n), .Q(
        StartOut) );
  DFFR_X2 done0_reg ( .D(\U3/U4/Z_0 ), .CK(clock), .RN(n622), .Q(n424) );
  DFFR_X2 \ReadAddress_reg[12]  ( .D(n712), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_12 ), .QN(n684) );
  DFFR_X2 \ReadAddress_reg[10]  ( .D(n714), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_10 ), .QN(n675) );
  DFFR_X2 \ReadAddress_reg[8]  ( .D(n716), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_8 ), .QN(n666) );
  DFFR_X2 \ReadAddress_reg[6]  ( .D(n718), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_6 ), .QN(n658) );
  DFFR_X2 \ReadAddress_reg[4]  ( .D(n720), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_4 ), .QN(n649) );
  DFFR_X2 \ReadAddress_reg[2]  ( .D(n722), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_2 ), .QN(n640) );
  DFFR_X2 \ReadAddress_reg[11]  ( .D(n713), .CK(clock), .RN(n627), .Q(
        \U4/DATA1_11 ), .QN(n632) );
  DFFR_X2 \ReadAddress_reg[9]  ( .D(n715), .CK(clock), .RN(n624), .Q(
        \U4/DATA1_9 ), .QN(n630) );
  DFFR_X2 \ReadAddress_reg[7]  ( .D(n717), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_7 ), .QN(n631) );
  DFFR_X2 \ReadAddress_reg[5]  ( .D(n719), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_5 ) );
  DFFR_X2 \ReadAddress_reg[3]  ( .D(n721), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_3 ) );
  DFFR_X2 \ReadAddress_reg[1]  ( .D(n723), .CK(clock), .RN(n623), .Q(
        \U4/DATA1_1 ) );
  DFFR_X2 \ReadAddress_reg[13]  ( .D(n711), .CK(clock), .RN(n622), .Q(
        \U4/DATA1_13 ), .QN(n688) );
  DFFR_X2 \ReadAddress_reg[14]  ( .D(n710), .CK(clock), .RN(n622), .Q(
        \U4/DATA1_14 ), .QN(n696) );
  INV_X4 U123 ( .A(1'b1), .ZN(DataOut[8]) );
  INV_X4 U125 ( .A(1'b1), .ZN(DataOut[9]) );
  INV_X4 U127 ( .A(1'b1), .ZN(DataOut[10]) );
  INV_X4 U129 ( .A(1'b1), .ZN(DataOut[11]) );
  INV_X4 U131 ( .A(1'b1), .ZN(DataOut[12]) );
  INV_X4 U133 ( .A(1'b1), .ZN(DataOut[13]) );
  INV_X4 U135 ( .A(1'b1), .ZN(DataOut[14]) );
  AND2_X4 U137 ( .A1(\U6/DATA1_1 ), .A2(n707), .ZN(n618) );
  OR2_X4 U138 ( .A1(n173), .A2(n174), .ZN(\U5/Z_7 ) );
  OR2_X4 U139 ( .A1(n199), .A2(n200), .ZN(\U5/Z_6 ) );
  OR2_X4 U140 ( .A1(n209), .A2(n210), .ZN(\U5/Z_5 ) );
  OR2_X4 U141 ( .A1(n219), .A2(n220), .ZN(\U5/Z_4 ) );
  OR2_X4 U142 ( .A1(n229), .A2(n230), .ZN(\U5/Z_3 ) );
  OR2_X4 U144 ( .A1(n239), .A2(n240), .ZN(\U5/Z_2 ) );
  OR2_X4 U145 ( .A1(n249), .A2(n250), .ZN(\U5/Z_1 ) );
  OR2_X4 U146 ( .A1(n259), .A2(n260), .ZN(\U5/Z_0 ) );
  NAND3_X1 U147 ( .A1(\U4/DATA1_1 ), .A2(\U4/DATA1_0 ), .A3(\U4/DATA1_2 ), 
        .ZN(n643) );
  INV_X4 U149 ( .A(n628), .ZN(n626) );
  INV_X4 U150 ( .A(n628), .ZN(n625) );
  INV_X4 U151 ( .A(n628), .ZN(n624) );
  INV_X4 U152 ( .A(n628), .ZN(n623) );
  INV_X4 U154 ( .A(n628), .ZN(n627) );
  INV_X4 U155 ( .A(n628), .ZN(n622) );
  INV_X4 U156 ( .A(reset_n), .ZN(n628) );
  OAI21_X2 U157 ( .B1(n708), .B2(n155), .A(n172), .ZN(\U3/U3/Z_0 ) );
  INV_X4 U159 ( .A(n621), .ZN(n619) );
  NAND2_X2 U160 ( .A1(n171), .A2(n635), .ZN(n693) );
  INV_X4 U161 ( .A(n629), .ZN(n709) );
  INV_X4 U162 ( .A(n621), .ZN(n620) );
  AOI21_X2 U164 ( .B1(n146), .B2(n726), .A(\U3/U4/Z_0 ), .ZN(n275) );
  OAI21_X2 U165 ( .B1(\U6/DATA1_1 ), .B2(n172), .A(n275), .ZN(n273) );
  OAI21_X2 U166 ( .B1(n149), .B2(n695), .A(n694), .ZN(n281) );
  OAI21_X2 U167 ( .B1(n727), .B2(n172), .A(n272), .ZN(\U3/U5/Z_3 ) );
  OAI21_X2 U169 ( .B1(n273), .B2(n726), .A(\U6/DATA1_3 ), .ZN(n272) );
  OAI21_X2 U170 ( .B1(n725), .B2(n707), .A(n274), .ZN(\U3/U5/Z_2 ) );
  OAI21_X2 U171 ( .B1(\U6/DATA1_0 ), .B2(n172), .A(n724), .ZN(\U3/U5/Z_0 ) );
  INV_X4 U172 ( .A(start), .ZN(n621) );
  AOI22_X2 U174 ( .A1(\U5/DATA6_0 ), .A2(n181), .B1(\U5/DATA5_0 ), .B2(n182), 
        .ZN(n263) );
  AOI22_X2 U175 ( .A1(\U5/DATA6_1 ), .A2(n181), .B1(\U5/DATA5_1 ), .B2(n182), 
        .ZN(n253) );
  AOI22_X2 U176 ( .A1(\U5/DATA6_2 ), .A2(n181), .B1(\U5/DATA5_2 ), .B2(n182), 
        .ZN(n243) );
  AOI22_X2 U177 ( .A1(\U5/DATA6_3 ), .A2(n181), .B1(\U5/DATA5_3 ), .B2(n182), 
        .ZN(n233) );
  AOI22_X2 U179 ( .A1(\U5/DATA6_4 ), .A2(n181), .B1(\U5/DATA5_4 ), .B2(n182), 
        .ZN(n223) );
  AOI22_X2 U180 ( .A1(\U5/DATA6_5 ), .A2(n181), .B1(\U5/DATA5_5 ), .B2(n182), 
        .ZN(n213) );
  AOI22_X2 U181 ( .A1(\U5/DATA6_6 ), .A2(n181), .B1(\U5/DATA5_6 ), .B2(n182), 
        .ZN(n203) );
  AOI22_X2 U182 ( .A1(\U5/DATA6_7 ), .A2(n181), .B1(\U5/DATA5_7 ), .B2(n182), 
        .ZN(n177) );
  AOI22_X2 U184 ( .A1(\U5/DATA10_0 ), .A2(n197), .B1(\U5/DATA9_0 ), .B2(n198), 
        .ZN(n268) );
  AOI22_X2 U185 ( .A1(\U5/DATA10_1 ), .A2(n197), .B1(\U5/DATA9_1 ), .B2(n198), 
        .ZN(n255) );
  AOI22_X2 U186 ( .A1(\U5/DATA10_2 ), .A2(n197), .B1(\U5/DATA9_2 ), .B2(n198), 
        .ZN(n245) );
  AOI22_X2 U187 ( .A1(\U5/DATA10_3 ), .A2(n197), .B1(\U5/DATA9_3 ), .B2(n198), 
        .ZN(n235) );
  AOI22_X2 U189 ( .A1(\U5/DATA10_4 ), .A2(n197), .B1(\U5/DATA9_4 ), .B2(n198), 
        .ZN(n225) );
  AOI22_X2 U190 ( .A1(\U5/DATA10_5 ), .A2(n197), .B1(\U5/DATA9_5 ), .B2(n198), 
        .ZN(n215) );
  AOI22_X2 U191 ( .A1(\U5/DATA10_6 ), .A2(n197), .B1(\U5/DATA9_6 ), .B2(n198), 
        .ZN(n205) );
  AOI22_X2 U192 ( .A1(\U5/DATA10_7 ), .A2(n197), .B1(\U5/DATA9_7 ), .B2(n198), 
        .ZN(n187) );
  AOI22_X2 U194 ( .A1(\U5/DATA2_0 ), .A2(n185), .B1(\U5/DATA1_0 ), .B2(n709), 
        .ZN(n261) );
  AOI22_X2 U195 ( .A1(\U5/DATA2_1 ), .A2(n185), .B1(\U5/DATA1_1 ), .B2(n709), 
        .ZN(n251) );
  AOI22_X2 U196 ( .A1(\U5/DATA2_2 ), .A2(n185), .B1(\U5/DATA1_2 ), .B2(n709), 
        .ZN(n241) );
  AOI22_X2 U197 ( .A1(\U5/DATA2_3 ), .A2(n185), .B1(\U5/DATA1_3 ), .B2(n709), 
        .ZN(n231) );
  AOI22_X2 U199 ( .A1(\U5/DATA2_4 ), .A2(n185), .B1(\U5/DATA1_4 ), .B2(n709), 
        .ZN(n221) );
  AOI22_X2 U200 ( .A1(\U5/DATA2_5 ), .A2(n185), .B1(\U5/DATA1_5 ), .B2(n709), 
        .ZN(n211) );
  AOI22_X2 U201 ( .A1(\U5/DATA2_6 ), .A2(n185), .B1(\U5/DATA1_6 ), .B2(n709), 
        .ZN(n201) );
  AOI22_X2 U202 ( .A1(\U5/DATA2_7 ), .A2(n185), .B1(\U5/DATA1_7 ), .B2(n709), 
        .ZN(n175) );
  AOI22_X2 U204 ( .A1(\U5/DATA12_0 ), .A2(n195), .B1(\U5/DATA11_0 ), .B2(n196), 
        .ZN(n269) );
  AOI22_X2 U205 ( .A1(\U5/DATA4_0 ), .A2(n183), .B1(\U5/DATA3_0 ), .B2(n184), 
        .ZN(n262) );
  AOI22_X2 U206 ( .A1(\U5/DATA12_1 ), .A2(n195), .B1(\U5/DATA11_1 ), .B2(n196), 
        .ZN(n256) );
  AOI22_X2 U207 ( .A1(\U5/DATA4_1 ), .A2(n183), .B1(\U5/DATA3_1 ), .B2(n184), 
        .ZN(n252) );
  AOI22_X2 U209 ( .A1(\U5/DATA12_2 ), .A2(n195), .B1(\U5/DATA11_2 ), .B2(n196), 
        .ZN(n246) );
  AOI22_X2 U210 ( .A1(\U5/DATA4_2 ), .A2(n183), .B1(\U5/DATA3_2 ), .B2(n184), 
        .ZN(n242) );
  AOI22_X2 U211 ( .A1(\U5/DATA12_3 ), .A2(n195), .B1(\U5/DATA11_3 ), .B2(n196), 
        .ZN(n236) );
  AOI22_X2 U212 ( .A1(\U5/DATA4_3 ), .A2(n183), .B1(\U5/DATA3_3 ), .B2(n184), 
        .ZN(n232) );
  AOI22_X2 U214 ( .A1(\U5/DATA12_4 ), .A2(n195), .B1(\U5/DATA11_4 ), .B2(n196), 
        .ZN(n226) );
  AOI22_X2 U217 ( .A1(\U5/DATA4_4 ), .A2(n183), .B1(\U5/DATA3_4 ), .B2(n184), 
        .ZN(n222) );
  AOI22_X2 U220 ( .A1(\U5/DATA12_5 ), .A2(n195), .B1(\U5/DATA11_5 ), .B2(n196), 
        .ZN(n216) );
  AOI22_X2 U223 ( .A1(\U5/DATA4_5 ), .A2(n183), .B1(\U5/DATA3_5 ), .B2(n184), 
        .ZN(n212) );
  AOI22_X2 U226 ( .A1(\U5/DATA12_6 ), .A2(n195), .B1(\U5/DATA11_6 ), .B2(n196), 
        .ZN(n206) );
  AOI22_X2 U229 ( .A1(\U5/DATA4_6 ), .A2(n183), .B1(\U5/DATA3_6 ), .B2(n184), 
        .ZN(n202) );
  AOI22_X2 U232 ( .A1(\U5/DATA12_7 ), .A2(n195), .B1(\U5/DATA11_7 ), .B2(n196), 
        .ZN(n188) );
  AOI22_X2 U235 ( .A1(\U5/DATA4_7 ), .A2(n183), .B1(\U5/DATA3_7 ), .B2(n184), 
        .ZN(n176) );
  AOI22_X2 U238 ( .A1(\U5/DATA16_0 ), .A2(n191), .B1(\U5/DATA15_0 ), .B2(n192), 
        .ZN(n271) );
  AOI22_X2 U239 ( .A1(\U5/DATA14_0 ), .A2(n193), .B1(\U5/DATA13_0 ), .B2(n194), 
        .ZN(n270) );
  AOI22_X2 U241 ( .A1(\U5/DATA8_0 ), .A2(n179), .B1(\U5/DATA7_0 ), .B2(n180), 
        .ZN(n264) );
  AOI22_X2 U242 ( .A1(\U5/DATA16_1 ), .A2(n191), .B1(\U5/DATA15_1 ), .B2(n192), 
        .ZN(n258) );
  AOI22_X2 U243 ( .A1(\U5/DATA14_1 ), .A2(n193), .B1(\U5/DATA13_1 ), .B2(n194), 
        .ZN(n257) );
  AOI22_X2 U244 ( .A1(\U5/DATA8_1 ), .A2(n179), .B1(\U5/DATA7_1 ), .B2(n180), 
        .ZN(n254) );
  AOI22_X2 U246 ( .A1(\U5/DATA16_2 ), .A2(n191), .B1(\U5/DATA15_2 ), .B2(n192), 
        .ZN(n248) );
  AOI22_X2 U248 ( .A1(\U5/DATA14_2 ), .A2(n193), .B1(\U5/DATA13_2 ), .B2(n194), 
        .ZN(n247) );
  AOI22_X2 U250 ( .A1(\U5/DATA8_2 ), .A2(n179), .B1(\U5/DATA7_2 ), .B2(n180), 
        .ZN(n244) );
  AOI22_X2 U251 ( .A1(\U5/DATA16_3 ), .A2(n191), .B1(\U5/DATA15_3 ), .B2(n192), 
        .ZN(n238) );
  AOI22_X2 U252 ( .A1(\U5/DATA14_3 ), .A2(n193), .B1(\U5/DATA13_3 ), .B2(n194), 
        .ZN(n237) );
  AOI22_X2 U253 ( .A1(\U5/DATA8_3 ), .A2(n179), .B1(\U5/DATA7_3 ), .B2(n180), 
        .ZN(n234) );
  AOI22_X2 U254 ( .A1(\U5/DATA16_4 ), .A2(n191), .B1(\U5/DATA15_4 ), .B2(n192), 
        .ZN(n228) );
  AOI22_X2 U255 ( .A1(\U5/DATA14_4 ), .A2(n193), .B1(\U5/DATA13_4 ), .B2(n194), 
        .ZN(n227) );
  AOI22_X2 U256 ( .A1(\U5/DATA8_4 ), .A2(n179), .B1(\U5/DATA7_4 ), .B2(n180), 
        .ZN(n224) );
  AOI22_X2 U257 ( .A1(\U5/DATA16_5 ), .A2(n191), .B1(\U5/DATA15_5 ), .B2(n192), 
        .ZN(n218) );
  AOI22_X2 U258 ( .A1(\U5/DATA14_5 ), .A2(n193), .B1(\U5/DATA13_5 ), .B2(n194), 
        .ZN(n217) );
  AOI22_X2 U259 ( .A1(\U5/DATA8_5 ), .A2(n179), .B1(\U5/DATA7_5 ), .B2(n180), 
        .ZN(n214) );
  AOI22_X2 U260 ( .A1(\U5/DATA16_6 ), .A2(n191), .B1(\U5/DATA15_6 ), .B2(n192), 
        .ZN(n208) );
  AOI22_X2 U261 ( .A1(\U5/DATA14_6 ), .A2(n193), .B1(\U5/DATA13_6 ), .B2(n194), 
        .ZN(n207) );
  AOI22_X2 U262 ( .A1(\U5/DATA8_6 ), .A2(n179), .B1(\U5/DATA7_6 ), .B2(n180), 
        .ZN(n204) );
  AOI22_X2 U263 ( .A1(\U5/DATA16_7 ), .A2(n191), .B1(\U5/DATA15_7 ), .B2(n192), 
        .ZN(n190) );
  AOI22_X2 U264 ( .A1(\U5/DATA14_7 ), .A2(n193), .B1(\U5/DATA13_7 ), .B2(n194), 
        .ZN(n189) );
  AOI22_X2 U265 ( .A1(\U5/DATA8_7 ), .A2(n179), .B1(\U5/DATA7_7 ), .B2(n180), 
        .ZN(n178) );
  NAND3_X1 U266 ( .A1(\U3/U2/DATA2_15 ), .A2(n155), .A3(n172), .ZN(n706) );
  NAND4_X2 U267 ( .A1(\U6/DATA1_2 ), .A2(\U6/DATA1_0 ), .A3(\U6/DATA1_3 ), 
        .A4(\U6/DATA1_1 ), .ZN(n629) );
  NAND2_X2 U268 ( .A1(n619), .A2(n629), .ZN(n172) );
  NAND2_X2 U269 ( .A1(n709), .A2(n619), .ZN(n155) );
  INV_X4 U270 ( .A(n643), .ZN(n646) );
  NAND3_X2 U271 ( .A1(\U4/DATA1_4 ), .A2(\U4/DATA1_3 ), .A3(n646), .ZN(n652)
         );
  INV_X4 U272 ( .A(n652), .ZN(n655) );
  NAND3_X2 U273 ( .A1(\U4/DATA1_6 ), .A2(\U4/DATA1_5 ), .A3(n655), .ZN(n661)
         );
  INV_X4 U274 ( .A(n661), .ZN(n669) );
  NOR3_X2 U275 ( .A1(n632), .A2(n631), .A3(n630), .ZN(n634) );
  NOR4_X2 U276 ( .A1(\U4/DATA1_10 ), .A2(\U4/DATA1_8 ), .A3(\U4/DATA1_13 ), 
        .A4(\U4/DATA1_12 ), .ZN(n633) );
  NAND4_X2 U277 ( .A1(\U4/DATA1_14 ), .A2(n669), .A3(n634), .A4(n633), .ZN(
        n171) );
  INV_X4 U278 ( .A(n155), .ZN(n635) );
  NOR2_X2 U279 ( .A1(n149), .A2(n693), .ZN(n637) );
  INV_X4 U280 ( .A(n171), .ZN(n708) );
  NAND2_X2 U281 ( .A1(n635), .A2(n708), .ZN(n636) );
  NAND2_X2 U282 ( .A1(n636), .A2(n172), .ZN(n698) );
  INV_X4 U283 ( .A(n698), .ZN(n695) );
  INV_X4 U284 ( .A(n693), .ZN(n702) );
  NAND2_X2 U285 ( .A1(n702), .A2(n149), .ZN(n694) );
  NAND2_X2 U286 ( .A1(n695), .A2(n694), .ZN(n639) );
  MUX2_X2 U287 ( .A(n637), .B(n639), .S(\U4/DATA1_1 ), .Z(n723) );
  NAND2_X2 U288 ( .A1(\U4/DATA1_0 ), .A2(n640), .ZN(n638) );
  MUX2_X2 U289 ( .A(n640), .B(n638), .S(\U4/DATA1_1 ), .Z(n642) );
  INV_X4 U290 ( .A(n639), .ZN(n641) );
  OAI22_X2 U291 ( .A1(n642), .A2(n693), .B1(n641), .B2(n640), .ZN(n722) );
  NOR2_X2 U292 ( .A1(n643), .A2(n693), .ZN(n645) );
  NAND2_X2 U293 ( .A1(n702), .A2(n643), .ZN(n644) );
  NAND2_X2 U294 ( .A1(n695), .A2(n644), .ZN(n648) );
  MUX2_X2 U295 ( .A(n645), .B(n648), .S(\U4/DATA1_3 ), .Z(n721) );
  NAND2_X2 U296 ( .A1(n646), .A2(n649), .ZN(n647) );
  MUX2_X2 U297 ( .A(n649), .B(n647), .S(\U4/DATA1_3 ), .Z(n651) );
  INV_X4 U298 ( .A(n648), .ZN(n650) );
  OAI22_X2 U299 ( .A1(n651), .A2(n693), .B1(n650), .B2(n649), .ZN(n720) );
  NOR2_X2 U300 ( .A1(n652), .A2(n693), .ZN(n654) );
  NAND2_X2 U301 ( .A1(n702), .A2(n652), .ZN(n653) );
  NAND2_X2 U302 ( .A1(n695), .A2(n653), .ZN(n657) );
  MUX2_X2 U303 ( .A(n654), .B(n657), .S(\U4/DATA1_5 ), .Z(n719) );
  NAND2_X2 U304 ( .A1(n655), .A2(n658), .ZN(n656) );
  MUX2_X2 U305 ( .A(n658), .B(n656), .S(\U4/DATA1_5 ), .Z(n660) );
  INV_X4 U306 ( .A(n657), .ZN(n659) );
  OAI22_X2 U307 ( .A1(n660), .A2(n693), .B1(n659), .B2(n658), .ZN(n718) );
  NOR2_X2 U308 ( .A1(n661), .A2(n693), .ZN(n663) );
  NAND2_X2 U309 ( .A1(n702), .A2(n661), .ZN(n662) );
  NAND2_X2 U310 ( .A1(n695), .A2(n662), .ZN(n665) );
  MUX2_X2 U311 ( .A(n663), .B(n665), .S(\U4/DATA1_7 ), .Z(n717) );
  NAND2_X2 U312 ( .A1(n669), .A2(n666), .ZN(n664) );
  MUX2_X2 U313 ( .A(n666), .B(n664), .S(\U4/DATA1_7 ), .Z(n668) );
  INV_X4 U314 ( .A(n665), .ZN(n667) );
  OAI22_X2 U315 ( .A1(n668), .A2(n693), .B1(n667), .B2(n666), .ZN(n716) );
  NAND3_X2 U316 ( .A1(\U4/DATA1_8 ), .A2(\U4/DATA1_7 ), .A3(n669), .ZN(n672)
         );
  NOR2_X2 U317 ( .A1(n672), .A2(n693), .ZN(n671) );
  NAND2_X2 U318 ( .A1(n702), .A2(n672), .ZN(n670) );
  NAND2_X2 U319 ( .A1(n695), .A2(n670), .ZN(n674) );
  MUX2_X2 U320 ( .A(n671), .B(n674), .S(\U4/DATA1_9 ), .Z(n715) );
  INV_X4 U321 ( .A(n672), .ZN(n678) );
  NAND2_X2 U322 ( .A1(n678), .A2(n675), .ZN(n673) );
  MUX2_X2 U323 ( .A(n675), .B(n673), .S(\U4/DATA1_9 ), .Z(n677) );
  INV_X4 U324 ( .A(n674), .ZN(n676) );
  OAI22_X2 U325 ( .A1(n677), .A2(n693), .B1(n676), .B2(n675), .ZN(n714) );
  NAND3_X2 U326 ( .A1(\U4/DATA1_10 ), .A2(\U4/DATA1_9 ), .A3(n678), .ZN(n681)
         );
  NOR2_X2 U327 ( .A1(n681), .A2(n693), .ZN(n680) );
  NAND2_X2 U328 ( .A1(n702), .A2(n681), .ZN(n679) );
  NAND2_X2 U329 ( .A1(n695), .A2(n679), .ZN(n683) );
  MUX2_X2 U330 ( .A(n680), .B(n683), .S(\U4/DATA1_11 ), .Z(n713) );
  INV_X4 U331 ( .A(n681), .ZN(n687) );
  NAND2_X2 U332 ( .A1(n687), .A2(n684), .ZN(n682) );
  MUX2_X2 U333 ( .A(n684), .B(n682), .S(\U4/DATA1_11 ), .Z(n686) );
  INV_X4 U334 ( .A(n683), .ZN(n685) );
  OAI22_X2 U335 ( .A1(n686), .A2(n693), .B1(n685), .B2(n684), .ZN(n712) );
  NAND3_X2 U336 ( .A1(\U4/DATA1_12 ), .A2(\U4/DATA1_11 ), .A3(n687), .ZN(n690)
         );
  XOR2_X2 U337 ( .A(n690), .B(\U4/DATA1_13 ), .Z(n689) );
  OAI22_X2 U338 ( .A1(n693), .A2(n689), .B1(n695), .B2(n688), .ZN(n711) );
  INV_X4 U339 ( .A(n690), .ZN(n691) );
  NAND2_X2 U340 ( .A1(\U4/DATA1_13 ), .A2(n691), .ZN(n700) );
  XOR2_X2 U341 ( .A(n700), .B(\U4/DATA1_14 ), .Z(n692) );
  OAI22_X2 U342 ( .A1(n693), .A2(n692), .B1(n695), .B2(n696), .ZN(n710) );
  NOR2_X2 U343 ( .A1(n696), .A2(n700), .ZN(n697) );
  NOR2_X2 U344 ( .A1(n155), .A2(n697), .ZN(n699) );
  NOR2_X2 U345 ( .A1(n699), .A2(n698), .ZN(n704) );
  INV_X4 U346 ( .A(n700), .ZN(n701) );
  NAND3_X2 U347 ( .A1(n702), .A2(\U4/DATA1_14 ), .A3(n701), .ZN(n703) );
  MUX2_X2 U348 ( .A(n704), .B(n703), .S(n147), .Z(n705) );
  NAND2_X2 U349 ( .A1(n706), .A2(n705), .ZN(n280) );
  NAND3_X2 U350 ( .A1(n726), .A2(\U6/DATA1_0 ), .A3(n618), .ZN(n274) );
  INV_X4 U351 ( .A(\U3/U4/Z_0 ), .ZN(n724) );
  INV_X4 U352 ( .A(n273), .ZN(n725) );
  INV_X4 U353 ( .A(n172), .ZN(n726) );
  INV_X4 U354 ( .A(n198), .ZN(n727) );
endmodule


module Output_Fetch_Cdf ( clock, reset_n, ReadBus, DataOut, StartIn, StartOut
 );
  input [127:0] ReadBus;
  output [19:0] DataOut;
  input clock, reset_n, StartIn;
  output StartOut;
  wire   \U3/U1/Z_0 ;
  assign \U3/U1/Z_0  = StartIn;

  DFF_X1 \DataOut_reg[19]  ( .D(ReadBus[19]), .CK(clock), .Q(DataOut[19]) );
  DFF_X1 \DataOut_reg[18]  ( .D(ReadBus[18]), .CK(clock), .Q(DataOut[18]) );
  DFF_X1 \DataOut_reg[17]  ( .D(ReadBus[17]), .CK(clock), .Q(DataOut[17]) );
  DFF_X1 \DataOut_reg[16]  ( .D(ReadBus[16]), .CK(clock), .Q(DataOut[16]) );
  DFF_X1 \DataOut_reg[15]  ( .D(ReadBus[15]), .CK(clock), .Q(DataOut[15]) );
  DFF_X1 \DataOut_reg[14]  ( .D(ReadBus[14]), .CK(clock), .Q(DataOut[14]) );
  DFF_X1 \DataOut_reg[13]  ( .D(ReadBus[13]), .CK(clock), .Q(DataOut[13]) );
  DFF_X1 \DataOut_reg[12]  ( .D(ReadBus[12]), .CK(clock), .Q(DataOut[12]) );
  DFF_X1 \DataOut_reg[11]  ( .D(ReadBus[11]), .CK(clock), .Q(DataOut[11]) );
  DFF_X1 \DataOut_reg[10]  ( .D(ReadBus[10]), .CK(clock), .Q(DataOut[10]) );
  DFF_X1 \DataOut_reg[9]  ( .D(ReadBus[9]), .CK(clock), .Q(DataOut[9]) );
  DFF_X1 \DataOut_reg[8]  ( .D(ReadBus[8]), .CK(clock), .Q(DataOut[8]) );
  DFF_X1 \DataOut_reg[7]  ( .D(ReadBus[7]), .CK(clock), .Q(DataOut[7]) );
  DFF_X1 \DataOut_reg[6]  ( .D(ReadBus[6]), .CK(clock), .Q(DataOut[6]) );
  DFF_X1 \DataOut_reg[5]  ( .D(ReadBus[5]), .CK(clock), .Q(DataOut[5]) );
  DFF_X1 \DataOut_reg[4]  ( .D(ReadBus[4]), .CK(clock), .Q(DataOut[4]) );
  DFF_X1 \DataOut_reg[3]  ( .D(ReadBus[3]), .CK(clock), .Q(DataOut[3]) );
  DFF_X1 \DataOut_reg[2]  ( .D(ReadBus[2]), .CK(clock), .Q(DataOut[2]) );
  DFF_X1 \DataOut_reg[1]  ( .D(ReadBus[1]), .CK(clock), .Q(DataOut[1]) );
  DFF_X1 \DataOut_reg[0]  ( .D(ReadBus[0]), .CK(clock), .Q(DataOut[0]) );
  DFFR_X2 StartOut_reg ( .D(\U3/U1/Z_0 ), .CK(clock), .RN(reset_n), .Q(
        StartOut) );
endmodule


module Output_TopExpression ( clock, reset_n, DataIn, CdfMin, StartIn, 
        StartOut, DataOut );
  input [19:0] DataIn;
  input [19:0] CdfMin;
  output [27:0] DataOut;
  input clock, reset_n, StartIn;
  output StartOut;
  wire   n81, n161, \U8/Z_0 , \U8/Z_1 , \U8/Z_2 , \U8/Z_3 , \U8/Z_4 , \U8/Z_5 ,
         \U8/Z_6 , \U8/Z_7 , \U8/Z_8 , \U8/Z_9 , \U8/Z_10 , \U8/Z_11 ,
         \U8/Z_12 , \U8/Z_13 , \U8/DATA1_8 , \U8/DATA1_9 , \U8/DATA1_10 ,
         \U8/DATA1_11 , \U8/DATA1_12 , \U8/DATA1_13 , \U7/Z_0 , \U7/Z_1 ,
         \U7/Z_2 , \U7/Z_3 , \U7/Z_4 , \U7/Z_5 , \U7/Z_6 , \U7/Z_7 , \U7/Z_8 ,
         \U7/Z_9 , \U7/Z_10 , \U7/Z_11 , \U7/Z_12 , \U7/Z_13 , \U7/Z_14 ,
         \U7/Z_15 , \U7/Z_16 , \U7/Z_17 , \U7/Z_19 , \U6/Z_0 , \U6/Z_1 ,
         \U6/Z_2 , \U6/Z_3 , \U6/Z_4 , \U6/Z_5 , \U6/Z_6 , \U6/Z_7 , \U6/Z_8 ,
         \U6/Z_9 , \U6/Z_10 , \U6/Z_11 , \U6/Z_12 , \U6/Z_13 , \U5/Z_0 ,
         \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 ,
         \U4/Z_7 , \U4/Z_8 , \U4/Z_9 , \U4/Z_10 , \U4/Z_11 , \U4/Z_12 ,
         \U4/Z_13 , \U4/Z_14 , \U4/Z_15 , \U4/Z_16 , \U4/Z_17 , \U4/Z_18 ,
         \U4/Z_19 , \U4/Z_20 , \U4/Z_21 , \U4/Z_22 , \U4/Z_23 , \U4/Z_24 ,
         \U4/Z_25 , \U4/Z_26 , \U4/Z_27 , \U4/DATA1_0 , \U4/DATA1_1 ,
         \U4/DATA1_2 , \U4/DATA1_3 , \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 ,
         \U4/DATA1_7 , \U4/DATA1_8 , \U4/DATA1_9 , \U4/DATA1_10 ,
         \U4/DATA1_11 , \U4/DATA1_12 , \U4/DATA1_13 , \top_add/CI ,
         \top_add/A[0] , \top_add/A[1] , \top_add/A[2] , \top_add/A[3] ,
         \top_add/A[4] , \top_add/A[5] , \top_add/A[11] , \top_add/A[12] ,
         \top_add/A[13] , \bottom_add/A[8] , \bottom_add/A[9] ,
         \bottom_add/A[10] , \bottom_add/A[11] , \bottom_add/A[12] ,
         \bottom_add/A[13] , \first_add/A[0] , \first_add/A[1] ,
         \first_add/A[2] , \first_add/A[3] , \first_add/A[4] ,
         \first_add/A[5] , \first_add/A[6] , \first_add/A[7] ,
         \first_add/A[8] , \first_add/A[9] , \first_add/A[10] ,
         \first_add/A[11] , \first_add/A[12] , \first_add/A[13] ,
         \first_add/A[14] , \first_add/A[15] , \first_add/A[16] ,
         \first_add/A[17] , \first_add/A[18] , \first_add/A[19] , n2, n3, n4,
         n5, n6, n7, n8, n9, n16, n17, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599;
  assign \first_add/A[0]  = DataIn[0];
  assign \first_add/A[1]  = DataIn[1];
  assign \first_add/A[2]  = DataIn[2];
  assign \first_add/A[3]  = DataIn[3];
  assign \first_add/A[4]  = DataIn[4];
  assign \first_add/A[5]  = DataIn[5];
  assign \first_add/A[6]  = DataIn[6];
  assign \first_add/A[7]  = DataIn[7];
  assign \first_add/A[8]  = DataIn[8];
  assign \first_add/A[9]  = DataIn[9];
  assign \first_add/A[10]  = DataIn[10];
  assign \first_add/A[11]  = DataIn[11];
  assign \first_add/A[12]  = DataIn[12];
  assign \first_add/A[13]  = DataIn[13];
  assign \first_add/A[14]  = DataIn[14];
  assign \first_add/A[15]  = DataIn[15];
  assign \first_add/A[16]  = DataIn[16];
  assign \first_add/A[17]  = DataIn[17];
  assign \first_add/A[18]  = DataIn[18];
  assign \first_add/A[19]  = DataIn[19];

  DFFR_X1 \Data_reg[19]  ( .D(\U7/Z_19 ), .CK(clock), .RN(n336), .Q(
        \U8/DATA1_13 ) );
  DFFR_X1 \DataOut_reg[26]  ( .D(\U4/Z_26 ), .CK(clock), .RN(n332), .Q(
        DataOut[26]) );
  AND2_X1 U75 ( .A1(\U4/DATA1_6 ), .A2(n81), .ZN(\U4/Z_6 ) );
  AND2_X1 U76 ( .A1(\U4/DATA1_5 ), .A2(n81), .ZN(\U4/Z_5 ) );
  AND2_X1 U77 ( .A1(\U4/DATA1_4 ), .A2(n81), .ZN(\U4/Z_4 ) );
  AND2_X1 U78 ( .A1(\U4/DATA1_3 ), .A2(n81), .ZN(\U4/Z_3 ) );
  AND2_X1 U87 ( .A1(\U4/DATA1_2 ), .A2(n81), .ZN(\U4/Z_2 ) );
  AND2_X1 U98 ( .A1(\U4/DATA1_1 ), .A2(n81), .ZN(\U4/Z_1 ) );
  AND2_X1 U99 ( .A1(\U4/DATA1_0 ), .A2(n81), .ZN(\U4/Z_0 ) );
  DFFR_X2 \dataTop_reg[19]  ( .D(\U8/Z_13 ), .CK(clock), .RN(n333), .Q(
        \top_add/A[13] ), .QN(n16) );
  DFFR_X2 \dataTop_reg[18]  ( .D(\U8/Z_12 ), .CK(clock), .RN(n333), .Q(
        \top_add/A[12] ), .QN(n17) );
  DFFR_X2 \dataTop_reg[17]  ( .D(\U8/Z_11 ), .CK(clock), .RN(n333), .Q(
        \top_add/A[11] ), .QN(n577) );
  DFFR_X2 \dataTop_reg[16]  ( .D(\U8/Z_10 ), .CK(clock), .RN(n333), .Q(n520), 
        .QN(n573) );
  DFFR_X2 \dataTop_reg[15]  ( .D(\U8/Z_9 ), .CK(clock), .RN(n333), .QN(n570)
         );
  DFFR_X2 \dataTop_reg[14]  ( .D(\U8/Z_8 ), .CK(clock), .RN(n333), .Q(n501), 
        .QN(n566) );
  DFFR_X2 \Data_reg[0]  ( .D(\U7/Z_0 ), .CK(clock), .RN(n334), .Q(
        \bottom_add/A[8] ), .QN(n412) );
  DFFR_X2 \Data_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .RN(n335), .Q(
        \bottom_add/A[9] ), .QN(n425) );
  DFFR_X2 \Data_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .RN(n335), .Q(
        \bottom_add/A[10] ), .QN(n441) );
  DFFR_X2 \Data_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .RN(n335), .Q(
        \bottom_add/A[11] ), .QN(n454) );
  DFFR_X2 \Data_reg[4]  ( .D(\U7/Z_4 ), .CK(clock), .RN(n335), .Q(
        \bottom_add/A[12] ), .QN(n470) );
  DFFR_X2 \Data_reg[5]  ( .D(\U7/Z_5 ), .CK(clock), .RN(n335), .Q(
        \bottom_add/A[13] ), .QN(n477) );
  DFFR_X2 \Data_reg[6]  ( .D(\U7/Z_6 ), .CK(clock), .RN(n335), .QN(n9) );
  DFFR_X2 \Data_reg[7]  ( .D(\U7/Z_7 ), .CK(clock), .RN(n335), .QN(n8) );
  DFFR_X2 \Data_reg[8]  ( .D(\U7/Z_8 ), .CK(clock), .RN(n335), .Q(n413), .QN(
        n7) );
  DFFR_X2 \Data_reg[9]  ( .D(\U7/Z_9 ), .CK(clock), .RN(n335), .Q(n426), .QN(
        n6) );
  DFFR_X2 \Data_reg[10]  ( .D(\U7/Z_10 ), .CK(clock), .RN(n335), .Q(n442), 
        .QN(n5) );
  DFFR_X2 \Data_reg[11]  ( .D(\U7/Z_11 ), .CK(clock), .RN(n335), .Q(n455), 
        .QN(n4) );
  DFFR_X2 \Data_reg[13]  ( .D(\U7/Z_13 ), .CK(clock), .RN(n336), .Q(n478), 
        .QN(n2) );
  DFFR_X2 \Data_reg[12]  ( .D(\U7/Z_12 ), .CK(clock), .RN(n335), .Q(n471), 
        .QN(n3) );
  DFFR_X2 Start0_reg ( .D(StartIn), .CK(clock), .RN(reset_n), .Q(n161), .QN(
        n598) );
  DFFR_X2 \dataTop_reg[7]  ( .D(\U8/Z_1 ), .CK(clock), .RN(n332), .Q(
        \top_add/A[1] ) );
  DFFR_X2 \dataTop_reg[6]  ( .D(\U8/Z_0 ), .CK(clock), .RN(n332), .Q(
        \top_add/A[0] ), .QN(n499) );
  DFFR_X2 \dataBottom_reg[0]  ( .D(\U6/Z_0 ), .CK(clock), .RN(n333), .Q(
        \U4/DATA1_0 ) );
  DFFR_X2 \dataTop_reg[13]  ( .D(\U8/Z_7 ), .CK(clock), .RN(n333), .QN(n563)
         );
  DFFR_X2 \dataTop_reg[12]  ( .D(\U8/Z_6 ), .CK(clock), .RN(n332), .QN(n560)
         );
  DFFR_X2 \dataTop_reg[11]  ( .D(\U8/Z_5 ), .CK(clock), .RN(n332), .Q(
        \top_add/A[5] ) );
  DFFR_X2 \dataTop_reg[10]  ( .D(\U8/Z_4 ), .CK(clock), .RN(n332), .Q(
        \top_add/A[4] ), .QN(n555) );
  DFFR_X2 \dataTop_reg[9]  ( .D(\U8/Z_3 ), .CK(clock), .RN(n332), .Q(
        \top_add/A[3] ) );
  DFFR_X2 \dataTop_reg[8]  ( .D(\U8/Z_2 ), .CK(clock), .RN(n332), .Q(
        \top_add/A[2] ), .QN(n519) );
  DFFR_X2 StartOut_reg ( .D(n81), .CK(clock), .RN(n332), .Q(StartOut) );
  DFFR_X2 \dataBottom_reg[1]  ( .D(\U6/Z_1 ), .CK(clock), .RN(n333), .Q(
        \U4/DATA1_1 ) );
  DFFR_X2 \DataOut_reg[13]  ( .D(\U4/Z_13 ), .CK(clock), .RN(n331), .Q(
        DataOut[13]) );
  DFFR_X2 \DataOut_reg[12]  ( .D(\U4/Z_12 ), .CK(clock), .RN(n331), .Q(
        DataOut[12]) );
  DFFR_X2 \DataOut_reg[11]  ( .D(\U4/Z_11 ), .CK(clock), .RN(reset_n), .Q(
        DataOut[11]) );
  DFFR_X2 \DataOut_reg[10]  ( .D(\U4/Z_10 ), .CK(clock), .RN(n336), .Q(
        DataOut[10]) );
  DFFR_X2 \DataOut_reg[9]  ( .D(\U4/Z_9 ), .CK(clock), .RN(n334), .Q(
        DataOut[9]) );
  DFFR_X2 \DataOut_reg[8]  ( .D(\U4/Z_8 ), .CK(clock), .RN(n335), .Q(
        DataOut[8]) );
  DFFR_X2 \DataOut_reg[7]  ( .D(\U4/Z_7 ), .CK(clock), .RN(n336), .Q(
        DataOut[7]) );
  DFFR_X2 \DataOut_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n334), .Q(
        DataOut[6]) );
  DFFR_X2 \DataOut_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n335), .Q(
        DataOut[5]) );
  DFFR_X2 \DataOut_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(n336), .Q(
        DataOut[4]) );
  DFFR_X2 \DataOut_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n336), .Q(
        DataOut[3]) );
  DFFR_X2 \DataOut_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .RN(n336), .Q(
        DataOut[2]) );
  DFFR_X2 \DataOut_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .RN(n336), .Q(
        DataOut[1]) );
  DFFR_X2 \DataOut_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n336), .Q(
        DataOut[0]) );
  DFFR_X2 \dataBottom_reg[2]  ( .D(\U6/Z_2 ), .CK(clock), .RN(n333), .Q(
        \U4/DATA1_2 ) );
  DFFR_X2 \dataBottom_reg[3]  ( .D(\U6/Z_3 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_3 ) );
  DFFR_X2 \dataBottom_reg[4]  ( .D(\U6/Z_4 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_4 ) );
  DFFR_X2 \dataBottom_reg[5]  ( .D(\U6/Z_5 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_5 ) );
  DFFR_X2 \DataOut_reg[15]  ( .D(\U4/Z_15 ), .CK(clock), .RN(n331), .Q(
        DataOut[15]) );
  DFFR_X2 \dataBottom_reg[6]  ( .D(\U6/Z_6 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_6 ) );
  DFFR_X2 \DataOut_reg[14]  ( .D(\U4/Z_14 ), .CK(clock), .RN(n331), .Q(
        DataOut[14]) );
  DFFR_X2 \dataBottom_reg[7]  ( .D(\U6/Z_7 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_7 ) );
  DFFR_X2 \dataBottom_reg[8]  ( .D(\U6/Z_8 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_8 ) );
  DFFR_X2 \DataOut_reg[16]  ( .D(\U4/Z_16 ), .CK(clock), .RN(n331), .Q(
        DataOut[16]) );
  DFFR_X2 \DataOut_reg[17]  ( .D(\U4/Z_17 ), .CK(clock), .RN(n331), .Q(
        DataOut[17]) );
  DFFR_X2 \dataBottom_reg[9]  ( .D(\U6/Z_9 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_9 ) );
  DFFR_X2 \dataBottom_reg[10]  ( .D(\U6/Z_10 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_10 ) );
  DFFR_X2 \DataOut_reg[18]  ( .D(\U4/Z_18 ), .CK(clock), .RN(n331), .Q(
        DataOut[18]) );
  DFFR_X2 \DataOut_reg[19]  ( .D(\U4/Z_19 ), .CK(clock), .RN(n331), .Q(
        DataOut[19]) );
  DFFR_X2 \dataBottom_reg[11]  ( .D(\U6/Z_11 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_11 ) );
  DFFR_X2 \DataOut_reg[20]  ( .D(\U4/Z_20 ), .CK(clock), .RN(n331), .Q(
        DataOut[20]) );
  DFFR_X2 \DataOut_reg[21]  ( .D(\U4/Z_21 ), .CK(clock), .RN(n331), .Q(
        DataOut[21]) );
  DFFR_X2 \dataBottom_reg[12]  ( .D(\U6/Z_12 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_12 ) );
  DFFR_X2 \Data_reg[14]  ( .D(\U7/Z_14 ), .CK(clock), .RN(n336), .Q(
        \U8/DATA1_8 ) );
  DFFR_X2 \Data_reg[15]  ( .D(\U7/Z_15 ), .CK(clock), .RN(n336), .Q(
        \U8/DATA1_9 ) );
  DFFR_X2 \DataOut_reg[25]  ( .D(\U4/Z_25 ), .CK(clock), .RN(n332), .Q(
        DataOut[25]) );
  DFFR_X2 \dataBottom_reg[13]  ( .D(\U6/Z_13 ), .CK(clock), .RN(n334), .Q(
        \U4/DATA1_13 ) );
  DFFR_X2 dataCout_reg ( .D(\U5/Z_0 ), .CK(clock), .RN(n333), .Q(\top_add/CI ), 
        .QN(n502) );
  DFFR_X2 Start1_reg ( .D(n161), .CK(clock), .RN(reset_n), .Q(n81), .QN(n584)
         );
  DFFR_X2 \DataOut_reg[22]  ( .D(\U4/Z_22 ), .CK(clock), .RN(n331), .Q(
        DataOut[22]) );
  DFFR_X2 \DataOut_reg[23]  ( .D(\U4/Z_23 ), .CK(clock), .RN(n331), .Q(
        DataOut[23]) );
  DFFR_X2 \DataOut_reg[24]  ( .D(\U4/Z_24 ), .CK(clock), .RN(n332), .Q(
        DataOut[24]) );
  DFFR_X2 \Data_reg[16]  ( .D(\U7/Z_16 ), .CK(clock), .RN(n336), .Q(
        \U8/DATA1_10 ) );
  DFFR_X2 \DataOut_reg[27]  ( .D(\U4/Z_27 ), .CK(clock), .RN(n332), .Q(
        DataOut[27]) );
  DFFR_X2 \Data_reg[17]  ( .D(\U7/Z_17 ), .CK(clock), .RN(n336), .Q(
        \U8/DATA1_11 ) );
  DFFR_X2 \Data_reg[18]  ( .D(n323), .CK(clock), .RN(n336), .Q(\U8/DATA1_12 )
         );
  NAND2_X1 U3 ( .A1(CdfMin[15]), .A2(n505), .ZN(n508) );
  INV_X1 U4 ( .A(CdfMin[17]), .ZN(n523) );
  NAND2_X2 U5 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X2 U6 ( .A1(n495), .A2(n496), .ZN(n507) );
  AOI22_X2 U7 ( .A1(n16), .A2(\top_add/A[5] ), .B1(n556), .B2(n308), .ZN(n322)
         );
  OAI21_X2 U8 ( .B1(\first_add/A[1] ), .B2(n342), .A(n384), .ZN(n343) );
  NOR2_X2 U9 ( .A1(\top_add/A[12] ), .A2(n582), .ZN(n583) );
  INV_X2 U10 ( .A(n521), .ZN(n534) );
  AOI22_X2 U11 ( .A1(n577), .A2(\top_add/A[3] ), .B1(n521), .B2(n305), .ZN(
        n321) );
  INV_X1 U12 ( .A(n503), .ZN(n511) );
  AOI22_X2 U13 ( .A1(n570), .A2(\top_add/A[1] ), .B1(n503), .B2(n304), .ZN(
        n320) );
  OR2_X4 U14 ( .A1(\top_add/A[1] ), .A2(n570), .ZN(n304) );
  OR2_X4 U15 ( .A1(\top_add/A[3] ), .A2(n577), .ZN(n305) );
  INV_X1 U16 ( .A(n556), .ZN(n559) );
  XNOR2_X2 U17 ( .A(n538), .B(CdfMin[18]), .ZN(n306) );
  INV_X4 U18 ( .A(CdfMin[1]), .ZN(n342) );
  AND2_X4 U19 ( .A1(n314), .A2(n566), .ZN(n307) );
  OAI221_X2 U20 ( .B1(\first_add/A[10] ), .B2(n436), .C1(n435), .C2(n434), .A(
        n433), .ZN(n459) );
  OR2_X4 U21 ( .A1(\top_add/A[5] ), .A2(n16), .ZN(n308) );
  AND2_X4 U22 ( .A1(n322), .A2(n560), .ZN(n315) );
  NOR2_X1 U23 ( .A1(n527), .A2(n526), .ZN(n533) );
  NAND2_X1 U24 ( .A1(n402), .A2(n401), .ZN(n392) );
  NOR2_X1 U25 ( .A1(n315), .A2(n561), .ZN(n562) );
  NAND2_X1 U26 ( .A1(\top_add/A[11] ), .A2(n579), .ZN(n580) );
  NOR2_X1 U27 ( .A1(n315), .A2(n563), .ZN(n564) );
  AND2_X2 U28 ( .A1(n315), .A2(n563), .ZN(n314) );
  XOR2_X1 U29 ( .A(n582), .B(\top_add/A[12] ), .Z(n581) );
  INV_X2 U30 ( .A(n359), .ZN(n355) );
  OAI221_X2 U31 ( .B1(\first_add/A[8] ), .B2(n407), .C1(n406), .C2(n405), .A(
        n404), .ZN(n430) );
  OAI221_X1 U32 ( .B1(\first_add/A[8] ), .B2(n407), .C1(n406), .C2(n405), .A(
        n404), .ZN(n309) );
  NAND3_X1 U33 ( .A1(n360), .A2(n359), .A3(n372), .ZN(n362) );
  NAND2_X2 U34 ( .A1(n508), .A2(n507), .ZN(n310) );
  NAND2_X2 U35 ( .A1(\first_add/A[15] ), .A2(n506), .ZN(n311) );
  AND2_X2 U36 ( .A1(n310), .A2(n311), .ZN(n514) );
  INV_X1 U37 ( .A(CdfMin[18]), .ZN(n536) );
  NAND2_X1 U38 ( .A1(n460), .A2(n459), .ZN(n447) );
  NAND2_X1 U39 ( .A1(CdfMin[17]), .A2(n524), .ZN(n529) );
  NAND2_X1 U40 ( .A1(CdfMin[2]), .A2(n380), .ZN(n345) );
  INV_X1 U41 ( .A(CdfMin[2]), .ZN(n340) );
  INV_X2 U42 ( .A(n525), .ZN(n528) );
  NAND2_X1 U43 ( .A1(n431), .A2(n309), .ZN(n418) );
  NAND2_X1 U44 ( .A1(n489), .A2(n488), .ZN(n481) );
  INV_X1 U45 ( .A(CdfMin[12]), .ZN(n465) );
  INV_X1 U46 ( .A(CdfMin[10]), .ZN(n436) );
  NOR2_X1 U47 ( .A1(CdfMin[0]), .A2(n386), .ZN(n387) );
  NAND2_X1 U48 ( .A1(CdfMin[18]), .A2(n538), .ZN(n549) );
  NAND2_X1 U49 ( .A1(CdfMin[6]), .A2(n347), .ZN(n349) );
  INV_X1 U50 ( .A(CdfMin[6]), .ZN(n338) );
  INV_X2 U51 ( .A(CdfMin[3]), .ZN(n341) );
  INV_X1 U52 ( .A(CdfMin[9]), .ZN(n419) );
  NAND2_X1 U53 ( .A1(CdfMin[9]), .A2(n417), .ZN(n433) );
  XNOR2_X1 U54 ( .A(CdfMin[9]), .B(\first_add/A[9] ), .ZN(n408) );
  INV_X1 U55 ( .A(CdfMin[14]), .ZN(n494) );
  INV_X1 U56 ( .A(CdfMin[15]), .ZN(n506) );
  XOR2_X2 U57 ( .A(n312), .B(n528), .Z(n517) );
  XOR2_X1 U58 ( .A(n524), .B(CdfMin[17]), .Z(n312) );
  XNOR2_X1 U59 ( .A(n497), .B(n507), .ZN(n498) );
  XOR2_X1 U60 ( .A(n505), .B(CdfMin[15]), .Z(n497) );
  XNOR2_X1 U61 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U62 ( .A(n380), .B(CdfMin[2]), .Z(n382) );
  XOR2_X1 U63 ( .A(n509), .B(n514), .Z(n510) );
  XNOR2_X1 U64 ( .A(CdfMin[16]), .B(\first_add/A[16] ), .ZN(n509) );
  XNOR2_X1 U65 ( .A(CdfMin[8]), .B(\first_add/A[8] ), .ZN(n316) );
  XNOR2_X1 U66 ( .A(CdfMin[10]), .B(\first_add/A[10] ), .ZN(n317) );
  XNOR2_X1 U67 ( .A(CdfMin[12]), .B(\first_add/A[12] ), .ZN(n318) );
  XNOR2_X1 U68 ( .A(CdfMin[14]), .B(\first_add/A[14] ), .ZN(n319) );
  XNOR2_X2 U69 ( .A(n313), .B(n388), .ZN(n385) );
  XOR2_X1 U70 ( .A(\first_add/A[1] ), .B(CdfMin[1]), .Z(n313) );
  XOR2_X1 U71 ( .A(\first_add/A[3] ), .B(CdfMin[3]), .Z(n324) );
  XOR2_X1 U72 ( .A(\first_add/A[5] ), .B(CdfMin[5]), .Z(n325) );
  XNOR2_X1 U73 ( .A(CdfMin[6]), .B(\first_add/A[6] ), .ZN(n326) );
  XNOR2_X1 U74 ( .A(n320), .B(n330), .ZN(n512) );
  XNOR2_X1 U79 ( .A(n534), .B(n327), .ZN(n522) );
  XNOR2_X1 U80 ( .A(n321), .B(n328), .ZN(n535) );
  XNOR2_X1 U81 ( .A(\top_add/A[1] ), .B(n570), .ZN(n329) );
  XNOR2_X1 U82 ( .A(n511), .B(n329), .ZN(n504) );
  INV_X4 U83 ( .A(n337), .ZN(n333) );
  INV_X4 U84 ( .A(n337), .ZN(n331) );
  INV_X4 U85 ( .A(n337), .ZN(n332) );
  INV_X4 U86 ( .A(n337), .ZN(n334) );
  INV_X4 U88 ( .A(n337), .ZN(n335) );
  INV_X4 U89 ( .A(n337), .ZN(n336) );
  INV_X4 U90 ( .A(reset_n), .ZN(n337) );
  AND2_X1 U91 ( .A1(n364), .A2(n361), .ZN(n352) );
  AND2_X1 U92 ( .A1(n515), .A2(CdfMin[16]), .ZN(n513) );
  AOI21_X1 U93 ( .B1(n582), .B2(n580), .A(n584), .ZN(\U4/Z_25 ) );
  XNOR2_X2 U94 ( .A(n395), .B(n316), .ZN(n396) );
  XNOR2_X2 U95 ( .A(n421), .B(n317), .ZN(n422) );
  XNOR2_X2 U96 ( .A(n450), .B(n318), .ZN(n451) );
  XNOR2_X2 U97 ( .A(n484), .B(n319), .ZN(n485) );
  AND4_X2 U100 ( .A1(n533), .A2(n532), .A3(n531), .A4(StartIn), .ZN(n323) );
  XOR2_X2 U101 ( .A(n324), .B(n378), .Z(n379) );
  XOR2_X2 U102 ( .A(n325), .B(n368), .Z(n369) );
  XNOR2_X2 U103 ( .A(n366), .B(n326), .ZN(n367) );
  XNOR2_X2 U104 ( .A(\top_add/A[3] ), .B(n577), .ZN(n327) );
  XNOR2_X2 U105 ( .A(\top_add/A[4] ), .B(n17), .ZN(n328) );
  INV_X4 U106 ( .A(StartIn), .ZN(n516) );
  XNOR2_X2 U107 ( .A(\top_add/A[2] ), .B(n573), .ZN(n330) );
  XNOR2_X2 U108 ( .A(CdfMin[7]), .B(\first_add/A[7] ), .ZN(n357) );
  NAND2_X2 U109 ( .A1(\first_add/A[6] ), .A2(n338), .ZN(n402) );
  INV_X4 U110 ( .A(\first_add/A[5] ), .ZN(n339) );
  NAND2_X2 U111 ( .A1(CdfMin[5]), .A2(n339), .ZN(n363) );
  NAND2_X2 U112 ( .A1(\first_add/A[2] ), .A2(n340), .ZN(n371) );
  NAND2_X2 U113 ( .A1(\first_add/A[3] ), .A2(n341), .ZN(n373) );
  INV_X4 U114 ( .A(\first_add/A[2] ), .ZN(n380) );
  NAND2_X2 U115 ( .A1(\first_add/A[1] ), .A2(n342), .ZN(n344) );
  INV_X4 U116 ( .A(\first_add/A[0] ), .ZN(n386) );
  NAND2_X2 U117 ( .A1(CdfMin[0]), .A2(n386), .ZN(n384) );
  NAND2_X2 U118 ( .A1(n344), .A2(n343), .ZN(n381) );
  NAND2_X2 U119 ( .A1(n345), .A2(n381), .ZN(n370) );
  NAND3_X2 U120 ( .A1(n371), .A2(n373), .A3(n370), .ZN(n359) );
  INV_X4 U121 ( .A(\first_add/A[4] ), .ZN(n346) );
  NAND2_X2 U122 ( .A1(CdfMin[4]), .A2(n346), .ZN(n360) );
  INV_X4 U123 ( .A(\first_add/A[6] ), .ZN(n347) );
  INV_X4 U124 ( .A(\first_add/A[3] ), .ZN(n348) );
  NAND2_X2 U125 ( .A1(CdfMin[3]), .A2(n348), .ZN(n372) );
  NAND3_X2 U126 ( .A1(n360), .A2(n349), .A3(n372), .ZN(n354) );
  INV_X4 U127 ( .A(n349), .ZN(n353) );
  INV_X4 U128 ( .A(CdfMin[5]), .ZN(n350) );
  NAND2_X2 U129 ( .A1(\first_add/A[5] ), .A2(n350), .ZN(n364) );
  INV_X4 U130 ( .A(CdfMin[4]), .ZN(n351) );
  NAND2_X2 U131 ( .A1(\first_add/A[4] ), .A2(n351), .ZN(n361) );
  OAI22_X2 U132 ( .A1(n355), .A2(n354), .B1(n353), .B2(n352), .ZN(n356) );
  NAND2_X2 U133 ( .A1(n356), .A2(n363), .ZN(n401) );
  XNOR2_X2 U134 ( .A(n357), .B(n392), .ZN(n358) );
  NOR2_X2 U135 ( .A1(n358), .A2(n516), .ZN(\U7/Z_7 ) );
  NAND2_X2 U136 ( .A1(n362), .A2(n361), .ZN(n368) );
  NAND2_X2 U137 ( .A1(n368), .A2(n363), .ZN(n365) );
  NAND2_X2 U138 ( .A1(n365), .A2(n364), .ZN(n366) );
  NOR2_X2 U139 ( .A1(n367), .A2(n516), .ZN(\U7/Z_6 ) );
  NOR2_X2 U140 ( .A1(n369), .A2(n516), .ZN(\U7/Z_5 ) );
  NAND2_X2 U141 ( .A1(n371), .A2(n370), .ZN(n378) );
  NAND2_X2 U142 ( .A1(n378), .A2(n372), .ZN(n374) );
  NAND2_X2 U143 ( .A1(n374), .A2(n373), .ZN(n376) );
  XOR2_X2 U144 ( .A(\first_add/A[4] ), .B(CdfMin[4]), .Z(n375) );
  XOR2_X2 U145 ( .A(n376), .B(n375), .Z(n377) );
  NOR2_X2 U146 ( .A1(n377), .A2(n516), .ZN(\U7/Z_4 ) );
  NOR2_X2 U147 ( .A1(n379), .A2(n516), .ZN(\U7/Z_3 ) );
  NOR2_X2 U148 ( .A1(n383), .A2(n516), .ZN(\U7/Z_2 ) );
  INV_X4 U149 ( .A(n384), .ZN(n388) );
  NOR2_X2 U150 ( .A1(n385), .A2(n516), .ZN(\U7/Z_1 ) );
  NOR2_X2 U151 ( .A1(n388), .A2(n387), .ZN(n389) );
  NOR2_X2 U152 ( .A1(n389), .A2(n516), .ZN(\U7/Z_0 ) );
  NAND3_X2 U153 ( .A1(n425), .A2(n441), .A3(n412), .ZN(n589) );
  INV_X4 U154 ( .A(n589), .ZN(n591) );
  NAND3_X2 U155 ( .A1(n454), .A2(n470), .A3(n591), .ZN(n594) );
  INV_X4 U156 ( .A(n594), .ZN(n596) );
  NAND3_X2 U157 ( .A1(n9), .A2(n477), .A3(n596), .ZN(n397) );
  XOR2_X2 U158 ( .A(n397), .B(n8), .Z(n390) );
  NOR2_X2 U159 ( .A1(n598), .A2(n390), .ZN(\U6/Z_7 ) );
  AND2_X1 U160 ( .A1(\U4/DATA1_7 ), .A2(n81), .ZN(\U4/Z_7 ) );
  INV_X4 U161 ( .A(\first_add/A[7] ), .ZN(n391) );
  NAND2_X2 U162 ( .A1(CdfMin[7]), .A2(n391), .ZN(n404) );
  NAND2_X2 U163 ( .A1(n392), .A2(n404), .ZN(n394) );
  INV_X4 U164 ( .A(CdfMin[7]), .ZN(n393) );
  NAND2_X2 U165 ( .A1(\first_add/A[7] ), .A2(n393), .ZN(n403) );
  NAND2_X2 U166 ( .A1(n394), .A2(n403), .ZN(n395) );
  NOR2_X2 U167 ( .A1(n396), .A2(n516), .ZN(\U7/Z_8 ) );
  XNOR2_X2 U168 ( .A(\bottom_add/A[8] ), .B(n7), .ZN(n399) );
  INV_X4 U169 ( .A(n397), .ZN(n398) );
  NAND2_X2 U170 ( .A1(n8), .A2(n398), .ZN(n410) );
  XNOR2_X2 U171 ( .A(n399), .B(n410), .ZN(n400) );
  NOR2_X2 U172 ( .A1(n400), .A2(n598), .ZN(\U6/Z_8 ) );
  AND2_X1 U173 ( .A1(\U4/DATA1_8 ), .A2(n81), .ZN(\U4/Z_8 ) );
  INV_X4 U174 ( .A(CdfMin[8]), .ZN(n407) );
  NAND2_X2 U175 ( .A1(\first_add/A[8] ), .A2(n407), .ZN(n431) );
  INV_X4 U176 ( .A(n401), .ZN(n406) );
  NAND2_X2 U177 ( .A1(n403), .A2(n402), .ZN(n405) );
  XNOR2_X2 U178 ( .A(n408), .B(n418), .ZN(n409) );
  NOR2_X2 U179 ( .A1(n409), .A2(n516), .ZN(\U7/Z_9 ) );
  NOR2_X2 U180 ( .A1(\bottom_add/A[8] ), .A2(n7), .ZN(n411) );
  OAI22_X2 U181 ( .A1(n413), .A2(n412), .B1(n411), .B2(n410), .ZN(n414) );
  INV_X4 U182 ( .A(n414), .ZN(n424) );
  XOR2_X2 U183 ( .A(\bottom_add/A[9] ), .B(n6), .Z(n415) );
  XOR2_X2 U184 ( .A(n424), .B(n415), .Z(n416) );
  NOR2_X2 U185 ( .A1(n416), .A2(n598), .ZN(\U6/Z_9 ) );
  AND2_X1 U186 ( .A1(\U4/DATA1_9 ), .A2(n81), .ZN(\U4/Z_9 ) );
  INV_X4 U187 ( .A(\first_add/A[9] ), .ZN(n417) );
  NAND2_X2 U188 ( .A1(n418), .A2(n433), .ZN(n420) );
  NAND2_X2 U189 ( .A1(\first_add/A[9] ), .A2(n419), .ZN(n432) );
  NAND2_X2 U190 ( .A1(n420), .A2(n432), .ZN(n421) );
  NOR2_X2 U191 ( .A1(n422), .A2(n516), .ZN(\U7/Z_10 ) );
  NOR2_X2 U192 ( .A1(\bottom_add/A[9] ), .A2(n6), .ZN(n423) );
  OAI22_X2 U193 ( .A1(n426), .A2(n425), .B1(n424), .B2(n423), .ZN(n427) );
  INV_X4 U194 ( .A(n427), .ZN(n440) );
  XOR2_X2 U195 ( .A(\bottom_add/A[10] ), .B(n5), .Z(n428) );
  XOR2_X2 U196 ( .A(n440), .B(n428), .Z(n429) );
  NOR2_X2 U197 ( .A1(n429), .A2(n598), .ZN(\U6/Z_10 ) );
  AND2_X1 U198 ( .A1(\U4/DATA1_10 ), .A2(n81), .ZN(\U4/Z_10 ) );
  XNOR2_X2 U199 ( .A(CdfMin[11]), .B(\first_add/A[11] ), .ZN(n437) );
  NAND2_X2 U200 ( .A1(\first_add/A[10] ), .A2(n436), .ZN(n460) );
  INV_X4 U201 ( .A(n430), .ZN(n435) );
  NAND2_X2 U202 ( .A1(n432), .A2(n431), .ZN(n434) );
  XNOR2_X2 U203 ( .A(n437), .B(n447), .ZN(n438) );
  NOR2_X2 U204 ( .A1(n438), .A2(n516), .ZN(\U7/Z_11 ) );
  NOR2_X2 U205 ( .A1(\bottom_add/A[10] ), .A2(n5), .ZN(n439) );
  OAI22_X2 U206 ( .A1(n442), .A2(n441), .B1(n440), .B2(n439), .ZN(n443) );
  INV_X4 U207 ( .A(n443), .ZN(n453) );
  XOR2_X2 U208 ( .A(\bottom_add/A[11] ), .B(n4), .Z(n444) );
  XOR2_X2 U209 ( .A(n453), .B(n444), .Z(n445) );
  NOR2_X2 U210 ( .A1(n445), .A2(n598), .ZN(\U6/Z_11 ) );
  AND2_X1 U211 ( .A1(\U4/DATA1_11 ), .A2(n81), .ZN(\U4/Z_11 ) );
  INV_X4 U212 ( .A(\first_add/A[11] ), .ZN(n446) );
  NAND2_X2 U213 ( .A1(CdfMin[11]), .A2(n446), .ZN(n462) );
  NAND2_X2 U214 ( .A1(n447), .A2(n462), .ZN(n449) );
  INV_X4 U215 ( .A(CdfMin[11]), .ZN(n448) );
  NAND2_X2 U216 ( .A1(\first_add/A[11] ), .A2(n448), .ZN(n461) );
  NAND2_X2 U217 ( .A1(n449), .A2(n461), .ZN(n450) );
  NOR2_X2 U218 ( .A1(n451), .A2(n516), .ZN(\U7/Z_12 ) );
  NOR2_X2 U219 ( .A1(\bottom_add/A[11] ), .A2(n4), .ZN(n452) );
  OAI22_X2 U220 ( .A1(n455), .A2(n454), .B1(n453), .B2(n452), .ZN(n456) );
  INV_X4 U221 ( .A(n456), .ZN(n469) );
  XOR2_X2 U222 ( .A(\bottom_add/A[12] ), .B(n3), .Z(n457) );
  XOR2_X2 U223 ( .A(n469), .B(n457), .Z(n458) );
  NOR2_X2 U224 ( .A1(n458), .A2(n598), .ZN(\U6/Z_12 ) );
  AND2_X1 U225 ( .A1(\U4/DATA1_12 ), .A2(n81), .ZN(\U4/Z_12 ) );
  XNOR2_X2 U226 ( .A(CdfMin[13]), .B(\first_add/A[13] ), .ZN(n466) );
  NAND2_X2 U227 ( .A1(\first_add/A[12] ), .A2(n465), .ZN(n489) );
  INV_X4 U228 ( .A(n459), .ZN(n464) );
  NAND2_X2 U229 ( .A1(n461), .A2(n460), .ZN(n463) );
  OAI221_X2 U230 ( .B1(\first_add/A[12] ), .B2(n465), .C1(n464), .C2(n463), 
        .A(n462), .ZN(n488) );
  XNOR2_X2 U231 ( .A(n466), .B(n481), .ZN(n467) );
  NOR2_X2 U232 ( .A1(n467), .A2(n516), .ZN(\U7/Z_13 ) );
  NOR2_X2 U233 ( .A1(\bottom_add/A[12] ), .A2(n3), .ZN(n468) );
  OAI22_X2 U234 ( .A1(n471), .A2(n470), .B1(n469), .B2(n468), .ZN(n472) );
  INV_X4 U235 ( .A(n472), .ZN(n476) );
  XOR2_X2 U236 ( .A(\bottom_add/A[13] ), .B(n2), .Z(n473) );
  XOR2_X2 U237 ( .A(n476), .B(n473), .Z(n474) );
  NOR2_X2 U238 ( .A1(n474), .A2(n598), .ZN(\U6/Z_13 ) );
  AND2_X1 U239 ( .A1(\U4/DATA1_13 ), .A2(n81), .ZN(\U4/Z_13 ) );
  NOR2_X2 U240 ( .A1(\bottom_add/A[13] ), .A2(n2), .ZN(n475) );
  OAI22_X2 U241 ( .A1(n478), .A2(n477), .B1(n476), .B2(n475), .ZN(n479) );
  AND2_X1 U242 ( .A1(n161), .A2(n479), .ZN(\U5/Z_0 ) );
  INV_X4 U243 ( .A(\first_add/A[13] ), .ZN(n480) );
  NAND2_X2 U244 ( .A1(CdfMin[13]), .A2(n480), .ZN(n491) );
  NAND2_X2 U245 ( .A1(n481), .A2(n491), .ZN(n483) );
  INV_X4 U246 ( .A(CdfMin[13]), .ZN(n482) );
  NAND2_X2 U247 ( .A1(\first_add/A[13] ), .A2(n482), .ZN(n490) );
  NAND2_X2 U248 ( .A1(n483), .A2(n490), .ZN(n484) );
  NOR2_X2 U249 ( .A1(n485), .A2(n516), .ZN(\U7/Z_14 ) );
  AND2_X1 U250 ( .A1(\U8/DATA1_8 ), .A2(n161), .ZN(\U8/Z_8 ) );
  NOR2_X2 U251 ( .A1(n598), .A2(n9), .ZN(\U8/Z_0 ) );
  XOR2_X2 U252 ( .A(n502), .B(n566), .Z(n486) );
  XOR2_X2 U253 ( .A(n486), .B(\top_add/A[0] ), .Z(n487) );
  NOR2_X2 U254 ( .A1(n487), .A2(n584), .ZN(\U4/Z_14 ) );
  NAND2_X2 U255 ( .A1(\first_add/A[14] ), .A2(n494), .ZN(n496) );
  INV_X4 U256 ( .A(n488), .ZN(n493) );
  NAND2_X2 U257 ( .A1(n490), .A2(n489), .ZN(n492) );
  OAI221_X2 U258 ( .B1(\first_add/A[14] ), .B2(n494), .C1(n493), .C2(n492), 
        .A(n491), .ZN(n495) );
  NOR2_X2 U259 ( .A1(n498), .A2(n516), .ZN(\U7/Z_15 ) );
  AND2_X1 U260 ( .A1(\U8/DATA1_9 ), .A2(n161), .ZN(\U8/Z_9 ) );
  NOR2_X2 U261 ( .A1(n598), .A2(n8), .ZN(\U8/Z_1 ) );
  NOR2_X2 U262 ( .A1(n566), .A2(\top_add/CI ), .ZN(n500) );
  OAI22_X2 U263 ( .A1(n502), .A2(n501), .B1(n500), .B2(n499), .ZN(n503) );
  NOR2_X2 U264 ( .A1(n504), .A2(n584), .ZN(\U4/Z_15 ) );
  INV_X4 U265 ( .A(\first_add/A[15] ), .ZN(n505) );
  NOR2_X2 U266 ( .A1(n510), .A2(n516), .ZN(\U7/Z_16 ) );
  AND2_X1 U267 ( .A1(\U8/DATA1_10 ), .A2(n161), .ZN(\U8/Z_10 ) );
  NOR2_X2 U268 ( .A1(n598), .A2(n7), .ZN(\U8/Z_2 ) );
  NOR2_X2 U269 ( .A1(n512), .A2(n584), .ZN(\U4/Z_16 ) );
  INV_X4 U270 ( .A(\first_add/A[17] ), .ZN(n524) );
  INV_X4 U271 ( .A(\first_add/A[16] ), .ZN(n515) );
  OAI22_X2 U272 ( .A1(CdfMin[16]), .A2(n515), .B1(n514), .B2(n513), .ZN(n525)
         );
  NOR2_X2 U273 ( .A1(n517), .A2(n516), .ZN(\U7/Z_17 ) );
  AND2_X1 U274 ( .A1(\U8/DATA1_11 ), .A2(n161), .ZN(\U8/Z_11 ) );
  NOR2_X2 U275 ( .A1(n598), .A2(n6), .ZN(\U8/Z_3 ) );
  NOR2_X2 U276 ( .A1(\top_add/A[2] ), .A2(n573), .ZN(n518) );
  OAI22_X2 U277 ( .A1(n520), .A2(n519), .B1(n320), .B2(n518), .ZN(n521) );
  NOR2_X2 U278 ( .A1(n522), .A2(n584), .ZN(\U4/Z_17 ) );
  INV_X4 U279 ( .A(\first_add/A[18] ), .ZN(n538) );
  NAND2_X2 U280 ( .A1(\first_add/A[17] ), .A2(n523), .ZN(n543) );
  NOR2_X2 U281 ( .A1(n306), .A2(n543), .ZN(n527) );
  NAND2_X2 U282 ( .A1(n525), .A2(n529), .ZN(n542) );
  NOR2_X2 U283 ( .A1(n306), .A2(n542), .ZN(n526) );
  NAND3_X2 U284 ( .A1(n543), .A2(n306), .A3(n528), .ZN(n532) );
  INV_X4 U285 ( .A(n529), .ZN(n530) );
  NAND2_X2 U286 ( .A1(n530), .A2(n306), .ZN(n531) );
  AND2_X1 U287 ( .A1(\U8/DATA1_12 ), .A2(n161), .ZN(\U8/Z_12 ) );
  NOR2_X2 U288 ( .A1(n598), .A2(n5), .ZN(\U8/Z_4 ) );
  NOR2_X2 U289 ( .A1(n535), .A2(n584), .ZN(\U4/Z_18 ) );
  NAND2_X2 U290 ( .A1(\first_add/A[18] ), .A2(n536), .ZN(n544) );
  INV_X4 U291 ( .A(n544), .ZN(n537) );
  XNOR2_X2 U292 ( .A(CdfMin[19]), .B(\first_add/A[19] ), .ZN(n548) );
  NAND2_X2 U293 ( .A1(n537), .A2(n548), .ZN(n541) );
  INV_X4 U294 ( .A(n549), .ZN(n539) );
  NAND2_X2 U295 ( .A1(n539), .A2(n545), .ZN(n540) );
  NAND3_X2 U296 ( .A1(n541), .A2(n540), .A3(StartIn), .ZN(n553) );
  NAND2_X2 U297 ( .A1(n543), .A2(n542), .ZN(n547) );
  INV_X4 U298 ( .A(n547), .ZN(n546) );
  INV_X4 U299 ( .A(n548), .ZN(n545) );
  NAND3_X2 U300 ( .A1(n546), .A2(n545), .A3(n544), .ZN(n551) );
  NAND3_X2 U301 ( .A1(n549), .A2(n548), .A3(n547), .ZN(n550) );
  NAND2_X2 U302 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X2 U303 ( .A1(n553), .A2(n552), .ZN(\U7/Z_19 ) );
  AND2_X1 U304 ( .A1(\U8/DATA1_13 ), .A2(n161), .ZN(\U8/Z_13 ) );
  NOR2_X2 U305 ( .A1(n598), .A2(n4), .ZN(\U8/Z_5 ) );
  NOR2_X2 U306 ( .A1(\top_add/A[4] ), .A2(n17), .ZN(n554) );
  OAI22_X2 U307 ( .A1(\top_add/A[12] ), .A2(n555), .B1(n321), .B2(n554), .ZN(
        n556) );
  XOR2_X2 U308 ( .A(\top_add/A[5] ), .B(n16), .Z(n557) );
  XOR2_X2 U309 ( .A(n559), .B(n557), .Z(n558) );
  NOR2_X2 U310 ( .A1(n558), .A2(n584), .ZN(\U4/Z_19 ) );
  NOR2_X2 U311 ( .A1(n598), .A2(n3), .ZN(\U8/Z_6 ) );
  NOR2_X2 U312 ( .A1(n322), .A2(n560), .ZN(n561) );
  NOR2_X2 U313 ( .A1(n562), .A2(n584), .ZN(\U4/Z_20 ) );
  NOR2_X2 U314 ( .A1(n598), .A2(n2), .ZN(\U8/Z_7 ) );
  NOR2_X2 U315 ( .A1(n314), .A2(n564), .ZN(n565) );
  NOR2_X2 U316 ( .A1(n565), .A2(n584), .ZN(\U4/Z_21 ) );
  NOR2_X2 U317 ( .A1(n314), .A2(n566), .ZN(n567) );
  NOR2_X2 U318 ( .A1(n307), .A2(n567), .ZN(n568) );
  NOR2_X2 U319 ( .A1(n568), .A2(n584), .ZN(\U4/Z_22 ) );
  NAND2_X2 U320 ( .A1(n307), .A2(n570), .ZN(n569) );
  INV_X4 U321 ( .A(n569), .ZN(n574) );
  NOR2_X2 U322 ( .A1(n307), .A2(n570), .ZN(n571) );
  NOR2_X2 U323 ( .A1(n574), .A2(n571), .ZN(n572) );
  NOR2_X2 U324 ( .A1(n572), .A2(n584), .ZN(\U4/Z_23 ) );
  NAND2_X2 U325 ( .A1(n574), .A2(n573), .ZN(n579) );
  INV_X4 U326 ( .A(n579), .ZN(n578) );
  NOR2_X2 U327 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X2 U328 ( .A1(n578), .A2(n575), .ZN(n576) );
  NOR2_X2 U329 ( .A1(n576), .A2(n584), .ZN(\U4/Z_24 ) );
  NOR2_X2 U330 ( .A1(n584), .A2(n581), .ZN(\U4/Z_26 ) );
  XNOR2_X2 U331 ( .A(n583), .B(\top_add/A[13] ), .ZN(n585) );
  NOR2_X2 U332 ( .A1(n585), .A2(n584), .ZN(\U4/Z_27 ) );
  NOR2_X2 U333 ( .A1(n598), .A2(n412), .ZN(\U6/Z_0 ) );
  XNOR2_X2 U334 ( .A(n425), .B(n412), .ZN(n586) );
  NOR2_X2 U335 ( .A1(n586), .A2(n598), .ZN(\U6/Z_1 ) );
  NAND2_X2 U336 ( .A1(n412), .A2(n425), .ZN(n587) );
  XOR2_X2 U337 ( .A(n587), .B(n441), .Z(n588) );
  NOR2_X2 U338 ( .A1(n598), .A2(n588), .ZN(\U6/Z_2 ) );
  XOR2_X2 U339 ( .A(n589), .B(n454), .Z(n590) );
  NOR2_X2 U340 ( .A1(n598), .A2(n590), .ZN(\U6/Z_3 ) );
  NAND2_X2 U341 ( .A1(n591), .A2(n454), .ZN(n592) );
  XOR2_X2 U342 ( .A(n592), .B(n470), .Z(n593) );
  NOR2_X2 U343 ( .A1(n598), .A2(n593), .ZN(\U6/Z_4 ) );
  XOR2_X2 U344 ( .A(n594), .B(n477), .Z(n595) );
  NOR2_X2 U345 ( .A1(n598), .A2(n595), .ZN(\U6/Z_5 ) );
  NAND2_X2 U346 ( .A1(n477), .A2(n596), .ZN(n597) );
  XOR2_X2 U347 ( .A(n597), .B(n9), .Z(n599) );
  NOR2_X2 U348 ( .A1(n599), .A2(n598), .ZN(\U6/Z_6 ) );
endmodule


module pipleline_stage_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n47, n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n87, n88, n89, n90, n91, n92, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n128, n129, n130, n131, n133, n134, n139, n141,
         n146, n147, n148, n150, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247;

  NAND2_X2 U4 ( .A1(n32), .A2(n25), .ZN(n23) );
  XNOR2_X2 U12 ( .A(n36), .B(n4), .ZN(SUM[18]) );
  XNOR2_X2 U28 ( .A(n43), .B(n6), .ZN(SUM[16]) );
  AOI21_X4 U29 ( .B1(n58), .B2(n39), .A(n40), .ZN(n1) );
  NAND2_X2 U32 ( .A1(n242), .A2(n42), .ZN(n6) );
  NAND2_X2 U35 ( .A1(B[16]), .A2(A[16]), .ZN(n42) );
  XNOR2_X2 U36 ( .A(n50), .B(n7), .ZN(SUM[15]) );
  NAND2_X2 U38 ( .A1(n226), .A2(n53), .ZN(n44) );
  NAND2_X2 U59 ( .A1(n66), .A2(n61), .ZN(n59) );
  AOI21_X4 U60 ( .B1(n218), .B2(n67), .A(n62), .ZN(n60) );
  NAND2_X2 U66 ( .A1(B[13]), .A2(A[13]), .ZN(n64) );
  XOR2_X2 U67 ( .A(n10), .B(n70), .Z(SUM[12]) );
  OAI21_X4 U70 ( .B1(n68), .B2(n74), .A(n69), .ZN(n67) );
  NAND2_X2 U71 ( .A1(n139), .A2(n69), .ZN(n10) );
  NAND2_X2 U74 ( .A1(B[12]), .A2(A[12]), .ZN(n69) );
  XNOR2_X2 U75 ( .A(n75), .B(n11), .ZN(SUM[11]) );
  NAND2_X2 U79 ( .A1(n71), .A2(n74), .ZN(n11) );
  NAND2_X2 U82 ( .A1(B[11]), .A2(A[11]), .ZN(n74) );
  XNOR2_X2 U83 ( .A(n81), .B(n12), .ZN(SUM[10]) );
  NAND2_X2 U88 ( .A1(n141), .A2(n80), .ZN(n12) );
  NOR2_X4 U90 ( .A1(B[10]), .A2(A[10]), .ZN(n79) );
  NAND2_X2 U91 ( .A1(B[10]), .A2(A[10]), .ZN(n80) );
  XNOR2_X2 U92 ( .A(n88), .B(n13), .ZN(SUM[9]) );
  XOR2_X2 U102 ( .A(n14), .B(n229), .Z(SUM[8]) );
  NAND2_X2 U111 ( .A1(B[8]), .A2(A[8]), .ZN(n90) );
  XOR2_X2 U112 ( .A(n15), .B(n103), .Z(SUM[7]) );
  OAI21_X4 U114 ( .B1(n114), .B2(n97), .A(n98), .ZN(n96) );
  NAND2_X2 U115 ( .A1(n104), .A2(n99), .ZN(n97) );
  NAND2_X2 U119 ( .A1(n99), .A2(n102), .ZN(n15) );
  XOR2_X2 U123 ( .A(n16), .B(n108), .Z(SUM[6]) );
  XNOR2_X2 U131 ( .A(n113), .B(n17), .ZN(SUM[5]) );
  NAND2_X2 U138 ( .A1(B[5]), .A2(A[5]), .ZN(n112) );
  XNOR2_X2 U139 ( .A(n119), .B(n18), .ZN(SUM[4]) );
  NAND2_X2 U144 ( .A1(n147), .A2(n118), .ZN(n18) );
  NAND2_X2 U147 ( .A1(B[4]), .A2(A[4]), .ZN(n118) );
  XOR2_X2 U148 ( .A(n19), .B(n122), .Z(SUM[3]) );
  NAND2_X2 U153 ( .A1(B[3]), .A2(A[3]), .ZN(n121) );
  NAND2_X2 U157 ( .A1(n234), .A2(n125), .ZN(n20) );
  NOR2_X4 U175 ( .A1(B[16]), .A2(A[16]), .ZN(n41) );
  XOR2_X1 U176 ( .A(n9), .B(n65), .Z(SUM[13]) );
  OAI21_X4 U177 ( .B1(n34), .B2(n38), .A(n35), .ZN(n219) );
  NOR2_X4 U178 ( .A1(B[18]), .A2(A[18]), .ZN(n34) );
  NAND2_X2 U179 ( .A1(n222), .A2(n107), .ZN(n105) );
  NAND2_X2 U180 ( .A1(n220), .A2(n221), .ZN(n222) );
  NAND2_X2 U181 ( .A1(B[14]), .A2(A[14]), .ZN(n52) );
  AOI21_X2 U182 ( .B1(n105), .B2(n99), .A(n100), .ZN(n98) );
  NAND2_X2 U183 ( .A1(n235), .A2(n125), .ZN(n123) );
  OAI21_X2 U184 ( .B1(n129), .B2(n131), .A(n130), .ZN(n224) );
  NOR2_X2 U185 ( .A1(n41), .A2(n44), .ZN(n39) );
  NAND2_X2 U186 ( .A1(B[7]), .A2(A[7]), .ZN(n102) );
  OR2_X4 U187 ( .A1(B[13]), .A2(A[13]), .ZN(n218) );
  OAI21_X1 U188 ( .B1(n34), .B2(n38), .A(n35), .ZN(n33) );
  INV_X2 U189 ( .A(n96), .ZN(n229) );
  NOR2_X2 U190 ( .A1(B[6]), .A2(A[6]), .ZN(n106) );
  NAND2_X1 U191 ( .A1(B[9]), .A2(A[9]), .ZN(n87) );
  INV_X1 U192 ( .A(n130), .ZN(n128) );
  NAND2_X2 U193 ( .A1(B[1]), .A2(A[1]), .ZN(n130) );
  NOR2_X2 U194 ( .A1(B[1]), .A2(A[1]), .ZN(n129) );
  NOR2_X2 U195 ( .A1(B[13]), .A2(A[13]), .ZN(n63) );
  INV_X4 U196 ( .A(n106), .ZN(n220) );
  INV_X4 U197 ( .A(n112), .ZN(n221) );
  NAND2_X1 U198 ( .A1(B[6]), .A2(A[6]), .ZN(n107) );
  INV_X1 U199 ( .A(n47), .ZN(n223) );
  INV_X2 U200 ( .A(n129), .ZN(n150) );
  INV_X1 U201 ( .A(n241), .ZN(n225) );
  OR2_X1 U202 ( .A1(A[15]), .A2(B[15]), .ZN(n226) );
  OR2_X1 U203 ( .A1(B[15]), .A2(A[15]), .ZN(n247) );
  OAI21_X2 U204 ( .B1(n1), .B2(n23), .A(n24), .ZN(CO) );
  INV_X4 U205 ( .A(n49), .ZN(n47) );
  NAND2_X4 U206 ( .A1(B[15]), .A2(A[15]), .ZN(n49) );
  NAND2_X1 U207 ( .A1(n146), .A2(n112), .ZN(n17) );
  NAND2_X1 U208 ( .A1(n91), .A2(n90), .ZN(n14) );
  INV_X4 U209 ( .A(n27), .ZN(n25) );
  NAND2_X1 U210 ( .A1(B[2]), .A2(A[2]), .ZN(n125) );
  AOI21_X1 U211 ( .B1(n150), .B2(n2), .A(n128), .ZN(n227) );
  INV_X1 U212 ( .A(n34), .ZN(n133) );
  OR2_X2 U213 ( .A1(B[9]), .A2(A[9]), .ZN(n246) );
  NAND2_X1 U214 ( .A1(n220), .A2(n107), .ZN(n16) );
  XNOR2_X1 U215 ( .A(n29), .B(n3), .ZN(SUM[19]) );
  OAI21_X2 U216 ( .B1(n245), .B2(n30), .A(n31), .ZN(n29) );
  AOI21_X2 U217 ( .B1(n219), .B2(n25), .A(n26), .ZN(n24) );
  INV_X1 U218 ( .A(n54), .ZN(n228) );
  NOR2_X2 U219 ( .A1(n34), .A2(n37), .ZN(n32) );
  INV_X2 U220 ( .A(n32), .ZN(n30) );
  INV_X4 U221 ( .A(n229), .ZN(n230) );
  NAND2_X2 U222 ( .A1(n237), .A2(n87), .ZN(n231) );
  INV_X4 U223 ( .A(n231), .ZN(n83) );
  NAND2_X2 U224 ( .A1(B[19]), .A2(A[19]), .ZN(n28) );
  AOI21_X4 U225 ( .B1(n96), .B2(n77), .A(n78), .ZN(n236) );
  OAI21_X1 U226 ( .B1(n106), .B2(n112), .A(n107), .ZN(n232) );
  OR2_X1 U227 ( .A1(B[9]), .A2(A[9]), .ZN(n233) );
  INV_X4 U228 ( .A(n90), .ZN(n92) );
  NOR2_X2 U229 ( .A1(B[3]), .A2(A[3]), .ZN(n120) );
  INV_X4 U230 ( .A(n63), .ZN(n61) );
  NAND2_X1 U231 ( .A1(n218), .A2(n64), .ZN(n9) );
  INV_X2 U232 ( .A(n64), .ZN(n62) );
  NAND2_X1 U233 ( .A1(n148), .A2(n121), .ZN(n19) );
  INV_X1 U234 ( .A(n120), .ZN(n148) );
  NAND2_X2 U235 ( .A1(B[17]), .A2(A[17]), .ZN(n38) );
  NAND2_X1 U236 ( .A1(n150), .A2(n130), .ZN(n21) );
  NAND2_X1 U237 ( .A1(n134), .A2(n38), .ZN(n5) );
  NAND2_X2 U238 ( .A1(n238), .A2(n239), .ZN(n240) );
  INV_X1 U239 ( .A(n37), .ZN(n134) );
  NOR2_X1 U240 ( .A1(B[17]), .A2(A[17]), .ZN(n37) );
  XOR2_X1 U241 ( .A(n8), .B(n57), .Z(SUM[14]) );
  NAND2_X2 U242 ( .A1(n224), .A2(n234), .ZN(n235) );
  INV_X4 U243 ( .A(n124), .ZN(n234) );
  INV_X1 U244 ( .A(n123), .ZN(n122) );
  NAND2_X2 U245 ( .A1(n243), .A2(n42), .ZN(n40) );
  INV_X1 U246 ( .A(n114), .ZN(n113) );
  NAND2_X1 U247 ( .A1(n233), .A2(n87), .ZN(n13) );
  NAND2_X1 U248 ( .A1(n233), .A2(n91), .ZN(n82) );
  AOI21_X4 U249 ( .B1(n247), .B2(n54), .A(n47), .ZN(n45) );
  OAI21_X4 U250 ( .B1(n121), .B2(n117), .A(n118), .ZN(n116) );
  AOI21_X1 U251 ( .B1(n230), .B2(n77), .A(n78), .ZN(n76) );
  OAI21_X4 U252 ( .B1(n83), .B2(n79), .A(n80), .ZN(n78) );
  NAND2_X2 U253 ( .A1(n246), .A2(n92), .ZN(n237) );
  INV_X1 U254 ( .A(n117), .ZN(n147) );
  NOR2_X4 U255 ( .A1(B[4]), .A2(A[4]), .ZN(n117) );
  NAND2_X4 U256 ( .A1(n240), .A2(n60), .ZN(n58) );
  INV_X4 U257 ( .A(n236), .ZN(n238) );
  INV_X4 U258 ( .A(n59), .ZN(n239) );
  INV_X1 U259 ( .A(n58), .ZN(n57) );
  AOI21_X4 U260 ( .B1(n123), .B2(n115), .A(n116), .ZN(n114) );
  INV_X2 U261 ( .A(n41), .ZN(n242) );
  INV_X4 U262 ( .A(n244), .ZN(n245) );
  NAND2_X2 U263 ( .A1(n241), .A2(n242), .ZN(n243) );
  INV_X4 U264 ( .A(n45), .ZN(n241) );
  AOI21_X1 U265 ( .B1(n113), .B2(n104), .A(n232), .ZN(n103) );
  AOI21_X1 U266 ( .B1(n75), .B2(n71), .A(n72), .ZN(n70) );
  INV_X1 U267 ( .A(n79), .ZN(n141) );
  INV_X1 U268 ( .A(n1), .ZN(n244) );
  AOI21_X1 U269 ( .B1(n75), .B2(n66), .A(n67), .ZN(n65) );
  NOR2_X2 U270 ( .A1(n82), .A2(n79), .ZN(n77) );
  NOR2_X2 U271 ( .A1(n117), .A2(n120), .ZN(n115) );
  AOI21_X2 U272 ( .B1(n113), .B2(n146), .A(n221), .ZN(n108) );
  OAI21_X1 U273 ( .B1(n122), .B2(n120), .A(n121), .ZN(n119) );
  OAI21_X1 U274 ( .B1(n229), .B2(n89), .A(n90), .ZN(n88) );
  OAI21_X1 U275 ( .B1(n229), .B2(n82), .A(n83), .ZN(n81) );
  NOR2_X2 U276 ( .A1(n68), .A2(n73), .ZN(n66) );
  NOR2_X2 U277 ( .A1(n106), .A2(n111), .ZN(n104) );
  NOR2_X2 U278 ( .A1(B[12]), .A2(A[12]), .ZN(n68) );
  NOR2_X1 U279 ( .A1(B[11]), .A2(A[11]), .ZN(n73) );
  NOR2_X1 U280 ( .A1(B[5]), .A2(A[5]), .ZN(n111) );
  NOR2_X1 U281 ( .A1(B[8]), .A2(A[8]), .ZN(n89) );
  NOR2_X2 U282 ( .A1(B[2]), .A2(A[2]), .ZN(n124) );
  NOR2_X2 U283 ( .A1(B[0]), .A2(A[0]), .ZN(n131) );
  NOR2_X2 U284 ( .A1(B[7]), .A2(A[7]), .ZN(n101) );
  NOR2_X2 U285 ( .A1(B[19]), .A2(A[19]), .ZN(n27) );
  OAI21_X1 U286 ( .B1(n57), .B2(n44), .A(n225), .ZN(n43) );
  NAND2_X1 U287 ( .A1(n226), .A2(n223), .ZN(n7) );
  NAND2_X1 U288 ( .A1(n25), .A2(n28), .ZN(n3) );
  NAND2_X1 U289 ( .A1(n133), .A2(n35), .ZN(n4) );
  NAND2_X2 U290 ( .A1(B[18]), .A2(A[18]), .ZN(n35) );
  NOR2_X1 U291 ( .A1(B[14]), .A2(A[14]), .ZN(n51) );
  XOR2_X1 U292 ( .A(n20), .B(n227), .Z(SUM[2]) );
  XOR2_X1 U293 ( .A(n131), .B(n21), .Z(SUM[1]) );
  XNOR2_X1 U294 ( .A(B[0]), .B(A[0]), .ZN(SUM[0]) );
  INV_X1 U295 ( .A(n33), .ZN(n31) );
  OAI21_X1 U296 ( .B1(n57), .B2(n51), .A(n228), .ZN(n50) );
  NAND2_X1 U297 ( .A1(n53), .A2(n228), .ZN(n8) );
  OAI21_X1 U298 ( .B1(n245), .B2(n37), .A(n38), .ZN(n36) );
  XOR2_X1 U299 ( .A(n5), .B(n245), .Z(SUM[17]) );
  INV_X4 U300 ( .A(n76), .ZN(n75) );
  INV_X4 U301 ( .A(n74), .ZN(n72) );
  INV_X4 U302 ( .A(n52), .ZN(n54) );
  INV_X4 U303 ( .A(n28), .ZN(n26) );
  INV_X4 U304 ( .A(n131), .ZN(n2) );
  INV_X4 U305 ( .A(n101), .ZN(n99) );
  INV_X4 U306 ( .A(n89), .ZN(n91) );
  INV_X4 U307 ( .A(n73), .ZN(n71) );
  INV_X4 U308 ( .A(n68), .ZN(n139) );
  INV_X4 U309 ( .A(n51), .ZN(n53) );
  INV_X4 U310 ( .A(n111), .ZN(n146) );
  INV_X4 U311 ( .A(n102), .ZN(n100) );
endmodule


module pipleline_stage_1 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151;
  wire   [20:0] stage_result;

  pipleline_stage_1_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(stage_out[0]) );
  INV_X4 U6 ( .A(n148), .ZN(q) );
  NAND2_X2 U7 ( .A1(divided[21]), .A2(n148), .ZN(n131) );
  NAND2_X2 U8 ( .A1(divided[22]), .A2(n126), .ZN(n129) );
  NAND2_X2 U9 ( .A1(divided[23]), .A2(n126), .ZN(n124) );
  NAND2_X2 U10 ( .A1(divided[24]), .A2(n148), .ZN(n120) );
  NAND2_X2 U11 ( .A1(divided[25]), .A2(n148), .ZN(n116) );
  NAND2_X2 U12 ( .A1(divided[13]), .A2(n126), .ZN(n127) );
  NAND2_X2 U13 ( .A1(divided[14]), .A2(n148), .ZN(n118) );
  NAND2_X2 U14 ( .A1(divided[15]), .A2(n107), .ZN(n122) );
  INV_X4 U15 ( .A(divided[27]), .ZN(n114) );
  INV_X4 U16 ( .A(n150), .ZN(n98) );
  INV_X4 U17 ( .A(n150), .ZN(n151) );
  INV_X1 U18 ( .A(n149), .ZN(n99) );
  INV_X4 U19 ( .A(n99), .ZN(n100) );
  NAND2_X2 U20 ( .A1(divided[11]), .A2(n126), .ZN(n101) );
  NAND2_X2 U21 ( .A1(stage_result[4]), .A2(q), .ZN(n102) );
  NAND2_X2 U22 ( .A1(n101), .A2(n102), .ZN(stage_out[12]) );
  NAND2_X2 U23 ( .A1(divided[10]), .A2(n148), .ZN(n103) );
  NAND2_X1 U24 ( .A1(stage_result[3]), .A2(q), .ZN(n104) );
  NAND2_X2 U25 ( .A1(n103), .A2(n104), .ZN(stage_out[11]) );
  NAND2_X2 U26 ( .A1(divided[12]), .A2(n126), .ZN(n105) );
  NAND2_X1 U27 ( .A1(stage_result[5]), .A2(q), .ZN(n106) );
  NAND2_X2 U28 ( .A1(n105), .A2(n106), .ZN(stage_out[13]) );
  NAND2_X2 U29 ( .A1(divided[18]), .A2(n107), .ZN(n108) );
  NAND2_X1 U30 ( .A1(stage_result[11]), .A2(q), .ZN(n109) );
  NAND2_X2 U31 ( .A1(n108), .A2(n109), .ZN(stage_out[19]) );
  INV_X1 U32 ( .A(q), .ZN(n107) );
  NAND2_X2 U33 ( .A1(divided[16]), .A2(n107), .ZN(n110) );
  NAND2_X1 U34 ( .A1(stage_result[9]), .A2(q), .ZN(n111) );
  NAND2_X2 U35 ( .A1(n110), .A2(n111), .ZN(stage_out[17]) );
  NAND2_X2 U36 ( .A1(divided[26]), .A2(n107), .ZN(n112) );
  NAND2_X1 U37 ( .A1(stage_result[19]), .A2(q), .ZN(n113) );
  NAND2_X2 U38 ( .A1(n112), .A2(n113), .ZN(stage_out[27]) );
  XNOR2_X2 U39 ( .A(n100), .B(n114), .ZN(n148) );
  XNOR2_X2 U40 ( .A(n149), .B(n114), .ZN(n150) );
  NAND2_X1 U41 ( .A1(stage_result[18]), .A2(q), .ZN(n117) );
  NAND2_X1 U42 ( .A1(n116), .A2(n117), .ZN(stage_out[26]) );
  NAND2_X1 U43 ( .A1(stage_result[7]), .A2(q), .ZN(n119) );
  NAND2_X1 U44 ( .A1(n118), .A2(n119), .ZN(stage_out[15]) );
  NAND2_X1 U45 ( .A1(stage_result[17]), .A2(q), .ZN(n121) );
  NAND2_X1 U46 ( .A1(n120), .A2(n121), .ZN(stage_out[25]) );
  NAND2_X1 U47 ( .A1(stage_result[8]), .A2(q), .ZN(n123) );
  NAND2_X1 U48 ( .A1(n122), .A2(n123), .ZN(stage_out[16]) );
  NAND2_X1 U49 ( .A1(stage_result[16]), .A2(q), .ZN(n125) );
  NAND2_X1 U50 ( .A1(n124), .A2(n125), .ZN(stage_out[24]) );
  NAND2_X1 U51 ( .A1(stage_result[6]), .A2(q), .ZN(n128) );
  NAND2_X1 U52 ( .A1(n127), .A2(n128), .ZN(stage_out[14]) );
  INV_X1 U53 ( .A(q), .ZN(n126) );
  NAND2_X1 U54 ( .A1(stage_result[15]), .A2(q), .ZN(n130) );
  NAND2_X1 U55 ( .A1(n129), .A2(n130), .ZN(stage_out[23]) );
  NAND2_X1 U56 ( .A1(stage_result[14]), .A2(q), .ZN(n132) );
  NAND2_X1 U57 ( .A1(n131), .A2(n132), .ZN(stage_out[22]) );
  NAND2_X1 U58 ( .A1(divided[17]), .A2(n148), .ZN(n142) );
  BUF_X4 U59 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U60 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U61 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U62 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U63 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U64 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U65 ( .A(divided[0]), .Z(stage_out[1]) );
  NAND2_X2 U66 ( .A1(divided[9]), .A2(n107), .ZN(n140) );
  NAND2_X1 U67 ( .A1(stage_result[2]), .A2(q), .ZN(n141) );
  NAND2_X1 U68 ( .A1(n140), .A2(n141), .ZN(stage_out[10]) );
  NAND2_X1 U69 ( .A1(stage_result[10]), .A2(q), .ZN(n143) );
  NAND2_X1 U70 ( .A1(n142), .A2(n143), .ZN(stage_out[18]) );
  NAND2_X2 U71 ( .A1(divided[8]), .A2(n148), .ZN(n144) );
  NAND2_X1 U72 ( .A1(stage_result[1]), .A2(q), .ZN(n145) );
  NAND2_X1 U73 ( .A1(n144), .A2(n145), .ZN(stage_out[9]) );
  NAND2_X2 U74 ( .A1(divided[7]), .A2(n148), .ZN(n146) );
  NAND2_X1 U75 ( .A1(stage_result[0]), .A2(q), .ZN(n147) );
  NAND2_X1 U76 ( .A1(n146), .A2(n147), .ZN(stage_out[8]) );
  INV_X4 U77 ( .A(stage_result[20]), .ZN(n149) );
  MUX2_X2 U78 ( .A(divided[19]), .B(stage_result[12]), .S(n151), .Z(
        stage_out[20]) );
  MUX2_X2 U79 ( .A(divided[20]), .B(stage_result[13]), .S(n98), .Z(
        stage_out[21]) );
endmodule


module pipleline_stage_7_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n38, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n129, n130, n131,
         n132, n133, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n211, n212, n213;

  XOR2_X2 U2 ( .A(n1), .B(n27), .Z(SUM[19]) );
  NAND2_X2 U4 ( .A1(n28), .A2(n212), .ZN(n21) );
  NAND2_X2 U8 ( .A1(n212), .A2(n26), .ZN(n1) );
  NAND2_X2 U11 ( .A1(A[19]), .A2(B[19]), .ZN(n26) );
  XOR2_X2 U12 ( .A(n2), .B(n32), .Z(SUM[18]) );
  NAND2_X2 U16 ( .A1(n126), .A2(n31), .ZN(n2) );
  NAND2_X2 U19 ( .A1(A[18]), .A2(B[18]), .ZN(n31) );
  XOR2_X2 U20 ( .A(n3), .B(n41), .Z(SUM[17]) );
  NAND2_X2 U24 ( .A1(n213), .A2(n211), .ZN(n35) );
  NAND2_X2 U28 ( .A1(n211), .A2(n40), .ZN(n3) );
  NAND2_X2 U31 ( .A1(A[17]), .A2(B[17]), .ZN(n40) );
  XNOR2_X2 U32 ( .A(n46), .B(n4), .ZN(SUM[16]) );
  NAND2_X2 U36 ( .A1(n213), .A2(n45), .ZN(n4) );
  NAND2_X2 U39 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U40 ( .A(n56), .B(n5), .ZN(SUM[15]) );
  NAND2_X2 U45 ( .A1(n60), .A2(n52), .ZN(n50) );
  NAND2_X2 U49 ( .A1(n129), .A2(n55), .ZN(n5) );
  NAND2_X2 U52 ( .A1(A[15]), .A2(B[15]), .ZN(n55) );
  XOR2_X2 U53 ( .A(n6), .B(n59), .Z(SUM[14]) );
  NAND2_X2 U55 ( .A1(n130), .A2(n58), .ZN(n6) );
  NAND2_X2 U58 ( .A1(A[14]), .A2(B[14]), .ZN(n58) );
  XNOR2_X2 U59 ( .A(n64), .B(n7), .ZN(SUM[13]) );
  NAND2_X2 U63 ( .A1(n131), .A2(n63), .ZN(n7) );
  NAND2_X2 U66 ( .A1(A[13]), .A2(B[13]), .ZN(n63) );
  XOR2_X2 U67 ( .A(n8), .B(n67), .Z(SUM[12]) );
  NAND2_X2 U69 ( .A1(n132), .A2(n66), .ZN(n8) );
  NAND2_X2 U72 ( .A1(A[12]), .A2(B[12]), .ZN(n66) );
  XOR2_X2 U73 ( .A(n9), .B(n75), .Z(SUM[11]) );
  NAND2_X2 U76 ( .A1(n83), .A2(n71), .ZN(n69) );
  NAND2_X2 U80 ( .A1(n133), .A2(n74), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[11]), .A2(B[11]), .ZN(n74) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[10]) );
  NAND2_X2 U88 ( .A1(n76), .A2(n79), .ZN(n10) );
  NAND2_X2 U91 ( .A1(A[10]), .A2(B[10]), .ZN(n79) );
  XNOR2_X2 U92 ( .A(n87), .B(n11), .ZN(SUM[9]) );
  NAND2_X2 U98 ( .A1(n135), .A2(n86), .ZN(n11) );
  NAND2_X2 U101 ( .A1(A[9]), .A2(B[9]), .ZN(n86) );
  XOR2_X2 U102 ( .A(n12), .B(n90), .Z(SUM[8]) );
  NAND2_X2 U104 ( .A1(n136), .A2(n89), .ZN(n12) );
  NAND2_X2 U107 ( .A1(A[8]), .A2(B[8]), .ZN(n89) );
  XNOR2_X2 U108 ( .A(n98), .B(n13), .ZN(SUM[7]) );
  NAND2_X2 U111 ( .A1(n102), .A2(n94), .ZN(n92) );
  NAND2_X2 U115 ( .A1(n137), .A2(n97), .ZN(n13) );
  NAND2_X2 U118 ( .A1(A[7]), .A2(B[7]), .ZN(n97) );
  XOR2_X2 U119 ( .A(n14), .B(n101), .Z(SUM[6]) );
  NAND2_X2 U121 ( .A1(n138), .A2(n100), .ZN(n14) );
  NAND2_X2 U124 ( .A1(A[6]), .A2(B[6]), .ZN(n100) );
  XOR2_X2 U125 ( .A(n15), .B(n106), .Z(SUM[5]) );
  NAND2_X2 U129 ( .A1(n139), .A2(n105), .ZN(n15) );
  NAND2_X2 U132 ( .A1(A[5]), .A2(B[5]), .ZN(n105) );
  XNOR2_X2 U133 ( .A(n111), .B(n16), .ZN(SUM[4]) );
  NAND2_X2 U137 ( .A1(n140), .A2(n110), .ZN(n16) );
  NAND2_X2 U140 ( .A1(A[4]), .A2(B[4]), .ZN(n110) );
  XNOR2_X2 U141 ( .A(n117), .B(n17), .ZN(SUM[3]) );
  NAND2_X2 U146 ( .A1(n141), .A2(n116), .ZN(n17) );
  NAND2_X2 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n116) );
  XOR2_X2 U150 ( .A(n18), .B(n120), .Z(SUM[2]) );
  NAND2_X2 U152 ( .A1(n142), .A2(n119), .ZN(n18) );
  NAND2_X2 U155 ( .A1(A[2]), .A2(B[2]), .ZN(n119) );
  XOR2_X2 U156 ( .A(n124), .B(n19), .Z(SUM[1]) );
  NAND2_X2 U159 ( .A1(n143), .A2(n123), .ZN(n19) );
  NAND2_X2 U162 ( .A1(A[1]), .A2(B[1]), .ZN(n123) );
  XNOR2_X2 U163 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U168 ( .B1(n68), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X2 U169 ( .B1(n91), .B2(n48), .A(n49), .ZN(n47) );
  NOR2_X2 U170 ( .A1(n69), .A2(n50), .ZN(n48) );
  OAI21_X2 U171 ( .B1(n70), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X2 U172 ( .B1(n90), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X2 U173 ( .B1(n46), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X2 U174 ( .B1(n46), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U175 ( .B1(n111), .B2(n102), .A(n103), .ZN(n101) );
  OAI21_X2 U176 ( .B1(n90), .B2(n81), .A(n82), .ZN(n80) );
  AOI21_X2 U177 ( .B1(n211), .B2(n43), .A(n38), .ZN(n36) );
  AOI21_X2 U178 ( .B1(n113), .B2(n121), .A(n114), .ZN(n112) );
  NOR2_X2 U179 ( .A1(n118), .A2(n115), .ZN(n113) );
  OAI21_X2 U180 ( .B1(n115), .B2(n119), .A(n116), .ZN(n114) );
  OAI21_X2 U181 ( .B1(n36), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X2 U182 ( .B1(n62), .B2(n66), .A(n63), .ZN(n61) );
  OAI21_X2 U183 ( .B1(n104), .B2(n110), .A(n105), .ZN(n103) );
  OAI21_X2 U184 ( .B1(n112), .B2(n92), .A(n93), .ZN(n91) );
  AOI21_X2 U185 ( .B1(n94), .B2(n103), .A(n95), .ZN(n93) );
  NOR2_X2 U186 ( .A1(n99), .A2(n96), .ZN(n94) );
  AOI21_X2 U187 ( .B1(n52), .B2(n61), .A(n53), .ZN(n51) );
  OAI21_X2 U188 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  AOI21_X2 U189 ( .B1(n29), .B2(n212), .A(n24), .ZN(n22) );
  AOI21_X2 U190 ( .B1(n46), .B2(n213), .A(n43), .ZN(n41) );
  OAI21_X2 U191 ( .B1(n122), .B2(n124), .A(n123), .ZN(n121) );
  OAI21_X2 U192 ( .B1(n85), .B2(n89), .A(n86), .ZN(n84) );
  OAI21_X2 U193 ( .B1(n96), .B2(n100), .A(n97), .ZN(n95) );
  AOI21_X2 U194 ( .B1(n71), .B2(n84), .A(n72), .ZN(n70) );
  OAI21_X2 U195 ( .B1(n73), .B2(n79), .A(n74), .ZN(n72) );
  OAI21_X2 U196 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X2 U197 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NOR2_X2 U198 ( .A1(n78), .A2(n73), .ZN(n71) );
  NOR2_X2 U199 ( .A1(n57), .A2(n54), .ZN(n52) );
  NOR2_X2 U200 ( .A1(n109), .A2(n104), .ZN(n102) );
  NOR2_X2 U201 ( .A1(n65), .A2(n62), .ZN(n60) );
  NOR2_X2 U202 ( .A1(n88), .A2(n85), .ZN(n83) );
  AOI21_X2 U203 ( .B1(n111), .B2(n140), .A(n108), .ZN(n106) );
  AOI21_X2 U204 ( .B1(n80), .B2(n76), .A(n77), .ZN(n75) );
  OAI21_X2 U205 ( .B1(n101), .B2(n99), .A(n100), .ZN(n98) );
  OAI21_X2 U206 ( .B1(n90), .B2(n88), .A(n89), .ZN(n87) );
  OAI21_X2 U207 ( .B1(n120), .B2(n118), .A(n119), .ZN(n117) );
  NOR2_X2 U208 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U209 ( .A1(A[3]), .A2(B[3]), .ZN(n115) );
  NOR2_X2 U210 ( .A1(A[7]), .A2(B[7]), .ZN(n96) );
  NOR2_X2 U211 ( .A1(A[5]), .A2(B[5]), .ZN(n104) );
  NOR2_X2 U212 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  NOR2_X2 U213 ( .A1(A[13]), .A2(B[13]), .ZN(n62) );
  NOR2_X2 U214 ( .A1(A[11]), .A2(B[11]), .ZN(n73) );
  NOR2_X2 U215 ( .A1(A[9]), .A2(B[9]), .ZN(n85) );
  NOR2_X2 U216 ( .A1(A[2]), .A2(B[2]), .ZN(n118) );
  NOR2_X2 U217 ( .A1(A[6]), .A2(B[6]), .ZN(n99) );
  NOR2_X2 U218 ( .A1(A[8]), .A2(B[8]), .ZN(n88) );
  NOR2_X2 U219 ( .A1(A[12]), .A2(B[12]), .ZN(n65) );
  NOR2_X2 U220 ( .A1(A[1]), .A2(B[1]), .ZN(n122) );
  NOR2_X2 U221 ( .A1(A[0]), .A2(B[0]), .ZN(n124) );
  NOR2_X2 U222 ( .A1(A[4]), .A2(B[4]), .ZN(n109) );
  NOR2_X2 U223 ( .A1(A[10]), .A2(B[10]), .ZN(n78) );
  OAI21_X2 U224 ( .B1(n47), .B2(n21), .A(n22), .ZN(CO) );
  OR2_X1 U225 ( .A1(A[17]), .A2(B[17]), .ZN(n211) );
  NOR2_X2 U226 ( .A1(A[18]), .A2(B[18]), .ZN(n30) );
  OR2_X1 U227 ( .A1(A[19]), .A2(B[19]), .ZN(n212) );
  OR2_X1 U228 ( .A1(A[16]), .A2(B[16]), .ZN(n213) );
  NOR2_X2 U229 ( .A1(A[14]), .A2(B[14]), .ZN(n57) );
  INV_X4 U230 ( .A(n91), .ZN(n90) );
  INV_X4 U231 ( .A(n84), .ZN(n82) );
  INV_X4 U232 ( .A(n83), .ZN(n81) );
  INV_X4 U233 ( .A(n79), .ZN(n77) );
  INV_X4 U234 ( .A(n68), .ZN(n67) );
  INV_X4 U235 ( .A(n47), .ZN(n46) );
  INV_X4 U236 ( .A(n45), .ZN(n43) );
  INV_X4 U237 ( .A(n40), .ZN(n38) );
  INV_X4 U238 ( .A(n36), .ZN(n34) );
  INV_X4 U239 ( .A(n35), .ZN(n33) );
  INV_X4 U240 ( .A(n26), .ZN(n24) );
  INV_X4 U241 ( .A(n122), .ZN(n143) );
  INV_X4 U242 ( .A(n118), .ZN(n142) );
  INV_X4 U243 ( .A(n115), .ZN(n141) );
  INV_X4 U244 ( .A(n104), .ZN(n139) );
  INV_X4 U245 ( .A(n99), .ZN(n138) );
  INV_X4 U246 ( .A(n96), .ZN(n137) );
  INV_X4 U247 ( .A(n88), .ZN(n136) );
  INV_X4 U248 ( .A(n85), .ZN(n135) );
  INV_X4 U249 ( .A(n78), .ZN(n76) );
  INV_X4 U250 ( .A(n73), .ZN(n133) );
  INV_X4 U251 ( .A(n65), .ZN(n132) );
  INV_X4 U252 ( .A(n62), .ZN(n131) );
  INV_X4 U253 ( .A(n57), .ZN(n130) );
  INV_X4 U254 ( .A(n54), .ZN(n129) );
  INV_X4 U255 ( .A(n30), .ZN(n126) );
  INV_X4 U256 ( .A(n121), .ZN(n120) );
  INV_X4 U257 ( .A(n112), .ZN(n111) );
  INV_X4 U258 ( .A(n110), .ZN(n108) );
  INV_X4 U259 ( .A(n109), .ZN(n140) );
endmodule


module pipleline_stage_7 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n105;
  wire   [20:0] stage_result;

  pipleline_stage_7_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(stage_out[0]) );
  INV_X4 U6 ( .A(n105), .ZN(q) );
  BUF_X4 U7 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U8 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U9 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U10 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U11 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U12 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U13 ( .A(divided[0]), .Z(stage_out[1]) );
  XNOR2_X2 U14 ( .A(divided[27]), .B(stage_result[20]), .ZN(n105) );
  MUX2_X2 U15 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U16 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U17 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U18 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U19 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U20 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U22 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U23 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U24 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U25 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U26 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U27 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U28 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U29 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U30 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U31 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U32 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U33 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U34 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_6_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n38, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n129, n130, n131,
         n132, n133, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n211, n212, n213;

  XOR2_X2 U2 ( .A(n1), .B(n27), .Z(SUM[19]) );
  NAND2_X2 U4 ( .A1(n28), .A2(n213), .ZN(n21) );
  NAND2_X2 U8 ( .A1(n213), .A2(n26), .ZN(n1) );
  NAND2_X2 U11 ( .A1(A[19]), .A2(B[19]), .ZN(n26) );
  XOR2_X2 U12 ( .A(n2), .B(n32), .Z(SUM[18]) );
  NAND2_X2 U16 ( .A1(n126), .A2(n31), .ZN(n2) );
  NAND2_X2 U19 ( .A1(A[18]), .A2(B[18]), .ZN(n31) );
  XOR2_X2 U20 ( .A(n3), .B(n41), .Z(SUM[17]) );
  NAND2_X2 U24 ( .A1(n212), .A2(n211), .ZN(n35) );
  NAND2_X2 U28 ( .A1(n211), .A2(n40), .ZN(n3) );
  NAND2_X2 U31 ( .A1(A[17]), .A2(B[17]), .ZN(n40) );
  XNOR2_X2 U32 ( .A(n46), .B(n4), .ZN(SUM[16]) );
  NAND2_X2 U36 ( .A1(n212), .A2(n45), .ZN(n4) );
  NAND2_X2 U39 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U40 ( .A(n56), .B(n5), .ZN(SUM[15]) );
  NAND2_X2 U45 ( .A1(n60), .A2(n52), .ZN(n50) );
  NAND2_X2 U49 ( .A1(n129), .A2(n55), .ZN(n5) );
  NAND2_X2 U52 ( .A1(A[15]), .A2(B[15]), .ZN(n55) );
  XOR2_X2 U53 ( .A(n6), .B(n59), .Z(SUM[14]) );
  NAND2_X2 U55 ( .A1(n130), .A2(n58), .ZN(n6) );
  NAND2_X2 U58 ( .A1(A[14]), .A2(B[14]), .ZN(n58) );
  XNOR2_X2 U59 ( .A(n64), .B(n7), .ZN(SUM[13]) );
  NAND2_X2 U63 ( .A1(n131), .A2(n63), .ZN(n7) );
  NAND2_X2 U66 ( .A1(A[13]), .A2(B[13]), .ZN(n63) );
  XOR2_X2 U67 ( .A(n8), .B(n67), .Z(SUM[12]) );
  NAND2_X2 U69 ( .A1(n132), .A2(n66), .ZN(n8) );
  NAND2_X2 U72 ( .A1(A[12]), .A2(B[12]), .ZN(n66) );
  XOR2_X2 U73 ( .A(n9), .B(n75), .Z(SUM[11]) );
  NAND2_X2 U76 ( .A1(n83), .A2(n71), .ZN(n69) );
  NAND2_X2 U80 ( .A1(n133), .A2(n74), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[11]), .A2(B[11]), .ZN(n74) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[10]) );
  NAND2_X2 U88 ( .A1(n76), .A2(n79), .ZN(n10) );
  NAND2_X2 U91 ( .A1(A[10]), .A2(B[10]), .ZN(n79) );
  XNOR2_X2 U92 ( .A(n87), .B(n11), .ZN(SUM[9]) );
  NAND2_X2 U98 ( .A1(n135), .A2(n86), .ZN(n11) );
  NAND2_X2 U101 ( .A1(A[9]), .A2(B[9]), .ZN(n86) );
  XOR2_X2 U102 ( .A(n12), .B(n90), .Z(SUM[8]) );
  NAND2_X2 U104 ( .A1(n136), .A2(n89), .ZN(n12) );
  NAND2_X2 U107 ( .A1(A[8]), .A2(B[8]), .ZN(n89) );
  XNOR2_X2 U108 ( .A(n98), .B(n13), .ZN(SUM[7]) );
  NAND2_X2 U111 ( .A1(n102), .A2(n94), .ZN(n92) );
  NAND2_X2 U115 ( .A1(n137), .A2(n97), .ZN(n13) );
  NAND2_X2 U118 ( .A1(A[7]), .A2(B[7]), .ZN(n97) );
  XOR2_X2 U119 ( .A(n14), .B(n101), .Z(SUM[6]) );
  NAND2_X2 U121 ( .A1(n138), .A2(n100), .ZN(n14) );
  NAND2_X2 U124 ( .A1(A[6]), .A2(B[6]), .ZN(n100) );
  XOR2_X2 U125 ( .A(n15), .B(n106), .Z(SUM[5]) );
  NAND2_X2 U129 ( .A1(n139), .A2(n105), .ZN(n15) );
  NAND2_X2 U132 ( .A1(A[5]), .A2(B[5]), .ZN(n105) );
  XNOR2_X2 U133 ( .A(n111), .B(n16), .ZN(SUM[4]) );
  NAND2_X2 U137 ( .A1(n140), .A2(n110), .ZN(n16) );
  NAND2_X2 U140 ( .A1(A[4]), .A2(B[4]), .ZN(n110) );
  XNOR2_X2 U141 ( .A(n117), .B(n17), .ZN(SUM[3]) );
  NAND2_X2 U146 ( .A1(n141), .A2(n116), .ZN(n17) );
  NAND2_X2 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n116) );
  XOR2_X2 U150 ( .A(n18), .B(n120), .Z(SUM[2]) );
  NAND2_X2 U152 ( .A1(n142), .A2(n119), .ZN(n18) );
  NAND2_X2 U155 ( .A1(A[2]), .A2(B[2]), .ZN(n119) );
  XOR2_X2 U156 ( .A(n124), .B(n19), .Z(SUM[1]) );
  NAND2_X2 U159 ( .A1(n143), .A2(n123), .ZN(n19) );
  NAND2_X2 U162 ( .A1(A[1]), .A2(B[1]), .ZN(n123) );
  XNOR2_X2 U163 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U168 ( .B1(n111), .B2(n102), .A(n103), .ZN(n101) );
  AOI21_X2 U169 ( .B1(n68), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X2 U170 ( .B1(n91), .B2(n48), .A(n49), .ZN(n47) );
  NOR2_X2 U171 ( .A1(n69), .A2(n50), .ZN(n48) );
  OAI21_X2 U172 ( .B1(n70), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X2 U173 ( .B1(n90), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U174 ( .B1(n90), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X2 U175 ( .B1(n46), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X2 U176 ( .B1(n46), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U177 ( .B1(n71), .B2(n84), .A(n72), .ZN(n70) );
  OAI21_X2 U178 ( .B1(n73), .B2(n79), .A(n74), .ZN(n72) );
  AOI21_X2 U179 ( .B1(n211), .B2(n43), .A(n38), .ZN(n36) );
  AOI21_X2 U180 ( .B1(n113), .B2(n121), .A(n114), .ZN(n112) );
  NOR2_X2 U181 ( .A1(n118), .A2(n115), .ZN(n113) );
  OAI21_X2 U182 ( .B1(n115), .B2(n119), .A(n116), .ZN(n114) );
  OAI21_X2 U183 ( .B1(n36), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X2 U184 ( .B1(n62), .B2(n66), .A(n63), .ZN(n61) );
  OAI21_X2 U185 ( .B1(n104), .B2(n110), .A(n105), .ZN(n103) );
  OAI21_X2 U186 ( .B1(n112), .B2(n92), .A(n93), .ZN(n91) );
  AOI21_X2 U187 ( .B1(n94), .B2(n103), .A(n95), .ZN(n93) );
  NOR2_X2 U188 ( .A1(n99), .A2(n96), .ZN(n94) );
  AOI21_X2 U189 ( .B1(n52), .B2(n61), .A(n53), .ZN(n51) );
  OAI21_X2 U190 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  AOI21_X2 U191 ( .B1(n29), .B2(n213), .A(n24), .ZN(n22) );
  AOI21_X2 U192 ( .B1(n80), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X2 U193 ( .B1(n46), .B2(n212), .A(n43), .ZN(n41) );
  OAI21_X2 U194 ( .B1(n122), .B2(n124), .A(n123), .ZN(n121) );
  OAI21_X2 U195 ( .B1(n85), .B2(n89), .A(n86), .ZN(n84) );
  OAI21_X2 U196 ( .B1(n96), .B2(n100), .A(n97), .ZN(n95) );
  OAI21_X2 U197 ( .B1(n101), .B2(n99), .A(n100), .ZN(n98) );
  OAI21_X2 U198 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X2 U199 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NOR2_X2 U200 ( .A1(n57), .A2(n54), .ZN(n52) );
  NOR2_X2 U201 ( .A1(n78), .A2(n73), .ZN(n71) );
  NOR2_X2 U202 ( .A1(n109), .A2(n104), .ZN(n102) );
  NOR2_X2 U203 ( .A1(n65), .A2(n62), .ZN(n60) );
  NOR2_X2 U204 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U205 ( .A1(n88), .A2(n85), .ZN(n83) );
  AOI21_X2 U206 ( .B1(n111), .B2(n140), .A(n108), .ZN(n106) );
  OAI21_X2 U207 ( .B1(n120), .B2(n118), .A(n119), .ZN(n117) );
  OAI21_X2 U208 ( .B1(n90), .B2(n88), .A(n89), .ZN(n87) );
  NOR2_X2 U209 ( .A1(A[3]), .A2(B[3]), .ZN(n115) );
  NOR2_X2 U210 ( .A1(A[7]), .A2(B[7]), .ZN(n96) );
  NOR2_X2 U211 ( .A1(A[5]), .A2(B[5]), .ZN(n104) );
  NOR2_X2 U212 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  NOR2_X2 U213 ( .A1(A[13]), .A2(B[13]), .ZN(n62) );
  NOR2_X2 U214 ( .A1(A[11]), .A2(B[11]), .ZN(n73) );
  NOR2_X2 U215 ( .A1(A[9]), .A2(B[9]), .ZN(n85) );
  NOR2_X2 U216 ( .A1(A[18]), .A2(B[18]), .ZN(n30) );
  NOR2_X2 U217 ( .A1(A[2]), .A2(B[2]), .ZN(n118) );
  NOR2_X2 U218 ( .A1(A[6]), .A2(B[6]), .ZN(n99) );
  NOR2_X2 U219 ( .A1(A[8]), .A2(B[8]), .ZN(n88) );
  NOR2_X2 U220 ( .A1(A[12]), .A2(B[12]), .ZN(n65) );
  NOR2_X2 U221 ( .A1(A[14]), .A2(B[14]), .ZN(n57) );
  NOR2_X2 U222 ( .A1(A[1]), .A2(B[1]), .ZN(n122) );
  NOR2_X2 U223 ( .A1(A[0]), .A2(B[0]), .ZN(n124) );
  NOR2_X2 U224 ( .A1(A[4]), .A2(B[4]), .ZN(n109) );
  NOR2_X2 U225 ( .A1(A[10]), .A2(B[10]), .ZN(n78) );
  OAI21_X2 U226 ( .B1(n47), .B2(n21), .A(n22), .ZN(CO) );
  OR2_X1 U227 ( .A1(A[17]), .A2(B[17]), .ZN(n211) );
  OR2_X1 U228 ( .A1(A[16]), .A2(B[16]), .ZN(n212) );
  OR2_X1 U229 ( .A1(A[19]), .A2(B[19]), .ZN(n213) );
  INV_X4 U230 ( .A(n91), .ZN(n90) );
  INV_X4 U231 ( .A(n84), .ZN(n82) );
  INV_X4 U232 ( .A(n83), .ZN(n81) );
  INV_X4 U233 ( .A(n79), .ZN(n77) );
  INV_X4 U234 ( .A(n68), .ZN(n67) );
  INV_X4 U235 ( .A(n47), .ZN(n46) );
  INV_X4 U236 ( .A(n45), .ZN(n43) );
  INV_X4 U237 ( .A(n40), .ZN(n38) );
  INV_X4 U238 ( .A(n36), .ZN(n34) );
  INV_X4 U239 ( .A(n35), .ZN(n33) );
  INV_X4 U240 ( .A(n26), .ZN(n24) );
  INV_X4 U241 ( .A(n122), .ZN(n143) );
  INV_X4 U242 ( .A(n118), .ZN(n142) );
  INV_X4 U243 ( .A(n115), .ZN(n141) );
  INV_X4 U244 ( .A(n104), .ZN(n139) );
  INV_X4 U245 ( .A(n99), .ZN(n138) );
  INV_X4 U246 ( .A(n96), .ZN(n137) );
  INV_X4 U247 ( .A(n88), .ZN(n136) );
  INV_X4 U248 ( .A(n85), .ZN(n135) );
  INV_X4 U249 ( .A(n78), .ZN(n76) );
  INV_X4 U250 ( .A(n73), .ZN(n133) );
  INV_X4 U251 ( .A(n65), .ZN(n132) );
  INV_X4 U252 ( .A(n62), .ZN(n131) );
  INV_X4 U253 ( .A(n57), .ZN(n130) );
  INV_X4 U254 ( .A(n54), .ZN(n129) );
  INV_X4 U255 ( .A(n30), .ZN(n126) );
  INV_X4 U256 ( .A(n121), .ZN(n120) );
  INV_X4 U257 ( .A(n112), .ZN(n111) );
  INV_X4 U258 ( .A(n110), .ZN(n108) );
  INV_X4 U259 ( .A(n109), .ZN(n140) );
endmodule


module pipleline_stage_6 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n105;
  wire   [20:0] stage_result;

  pipleline_stage_6_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(stage_out[0]) );
  INV_X4 U6 ( .A(n105), .ZN(q) );
  BUF_X4 U7 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U8 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U9 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U10 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U11 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U12 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U13 ( .A(divided[0]), .Z(stage_out[1]) );
  XNOR2_X2 U14 ( .A(divided[27]), .B(stage_result[20]), .ZN(n105) );
  MUX2_X2 U15 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U16 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U17 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U18 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U19 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U20 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U22 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U23 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U24 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U25 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U26 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U27 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U28 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U29 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U30 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U31 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U32 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U33 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U34 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n38, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n129, n130, n131,
         n132, n133, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n211, n212, n213;

  XOR2_X2 U2 ( .A(n1), .B(n27), .Z(SUM[19]) );
  NAND2_X2 U4 ( .A1(n28), .A2(n213), .ZN(n21) );
  NAND2_X2 U8 ( .A1(n213), .A2(n26), .ZN(n1) );
  NAND2_X2 U11 ( .A1(A[19]), .A2(B[19]), .ZN(n26) );
  XOR2_X2 U12 ( .A(n2), .B(n32), .Z(SUM[18]) );
  NAND2_X2 U16 ( .A1(n126), .A2(n31), .ZN(n2) );
  NAND2_X2 U19 ( .A1(A[18]), .A2(B[18]), .ZN(n31) );
  XOR2_X2 U20 ( .A(n3), .B(n41), .Z(SUM[17]) );
  NAND2_X2 U24 ( .A1(n212), .A2(n211), .ZN(n35) );
  NAND2_X2 U28 ( .A1(n211), .A2(n40), .ZN(n3) );
  NAND2_X2 U31 ( .A1(A[17]), .A2(B[17]), .ZN(n40) );
  XNOR2_X2 U32 ( .A(n46), .B(n4), .ZN(SUM[16]) );
  NAND2_X2 U36 ( .A1(n212), .A2(n45), .ZN(n4) );
  NAND2_X2 U39 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U40 ( .A(n56), .B(n5), .ZN(SUM[15]) );
  NAND2_X2 U45 ( .A1(n60), .A2(n52), .ZN(n50) );
  NAND2_X2 U49 ( .A1(n129), .A2(n55), .ZN(n5) );
  NAND2_X2 U52 ( .A1(A[15]), .A2(B[15]), .ZN(n55) );
  XOR2_X2 U53 ( .A(n6), .B(n59), .Z(SUM[14]) );
  NAND2_X2 U55 ( .A1(n130), .A2(n58), .ZN(n6) );
  NAND2_X2 U58 ( .A1(A[14]), .A2(B[14]), .ZN(n58) );
  XNOR2_X2 U59 ( .A(n64), .B(n7), .ZN(SUM[13]) );
  NAND2_X2 U63 ( .A1(n131), .A2(n63), .ZN(n7) );
  NAND2_X2 U66 ( .A1(A[13]), .A2(B[13]), .ZN(n63) );
  XOR2_X2 U67 ( .A(n8), .B(n67), .Z(SUM[12]) );
  NAND2_X2 U69 ( .A1(n132), .A2(n66), .ZN(n8) );
  NAND2_X2 U72 ( .A1(A[12]), .A2(B[12]), .ZN(n66) );
  XOR2_X2 U73 ( .A(n9), .B(n75), .Z(SUM[11]) );
  NAND2_X2 U76 ( .A1(n83), .A2(n71), .ZN(n69) );
  NAND2_X2 U80 ( .A1(n133), .A2(n74), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[11]), .A2(B[11]), .ZN(n74) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[10]) );
  NAND2_X2 U88 ( .A1(n76), .A2(n79), .ZN(n10) );
  NAND2_X2 U91 ( .A1(A[10]), .A2(B[10]), .ZN(n79) );
  XNOR2_X2 U92 ( .A(n87), .B(n11), .ZN(SUM[9]) );
  NAND2_X2 U98 ( .A1(n135), .A2(n86), .ZN(n11) );
  NAND2_X2 U101 ( .A1(A[9]), .A2(B[9]), .ZN(n86) );
  XOR2_X2 U102 ( .A(n12), .B(n90), .Z(SUM[8]) );
  NAND2_X2 U104 ( .A1(n136), .A2(n89), .ZN(n12) );
  NAND2_X2 U107 ( .A1(A[8]), .A2(B[8]), .ZN(n89) );
  XNOR2_X2 U108 ( .A(n98), .B(n13), .ZN(SUM[7]) );
  NAND2_X2 U111 ( .A1(n102), .A2(n94), .ZN(n92) );
  NAND2_X2 U115 ( .A1(n137), .A2(n97), .ZN(n13) );
  NAND2_X2 U118 ( .A1(A[7]), .A2(B[7]), .ZN(n97) );
  XOR2_X2 U119 ( .A(n14), .B(n101), .Z(SUM[6]) );
  NAND2_X2 U121 ( .A1(n138), .A2(n100), .ZN(n14) );
  NAND2_X2 U124 ( .A1(A[6]), .A2(B[6]), .ZN(n100) );
  XOR2_X2 U125 ( .A(n15), .B(n106), .Z(SUM[5]) );
  NAND2_X2 U129 ( .A1(n139), .A2(n105), .ZN(n15) );
  NAND2_X2 U132 ( .A1(A[5]), .A2(B[5]), .ZN(n105) );
  XNOR2_X2 U133 ( .A(n111), .B(n16), .ZN(SUM[4]) );
  NAND2_X2 U137 ( .A1(n140), .A2(n110), .ZN(n16) );
  NAND2_X2 U140 ( .A1(A[4]), .A2(B[4]), .ZN(n110) );
  XNOR2_X2 U141 ( .A(n117), .B(n17), .ZN(SUM[3]) );
  NAND2_X2 U146 ( .A1(n141), .A2(n116), .ZN(n17) );
  NAND2_X2 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n116) );
  XOR2_X2 U150 ( .A(n18), .B(n120), .Z(SUM[2]) );
  NAND2_X2 U152 ( .A1(n142), .A2(n119), .ZN(n18) );
  NAND2_X2 U155 ( .A1(A[2]), .A2(B[2]), .ZN(n119) );
  XOR2_X2 U156 ( .A(n124), .B(n19), .Z(SUM[1]) );
  NAND2_X2 U159 ( .A1(n143), .A2(n123), .ZN(n19) );
  NAND2_X2 U162 ( .A1(A[1]), .A2(B[1]), .ZN(n123) );
  XNOR2_X2 U163 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U168 ( .B1(n111), .B2(n102), .A(n103), .ZN(n101) );
  AOI21_X2 U169 ( .B1(n68), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X2 U170 ( .B1(n91), .B2(n48), .A(n49), .ZN(n47) );
  NOR2_X2 U171 ( .A1(n69), .A2(n50), .ZN(n48) );
  OAI21_X2 U172 ( .B1(n70), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X2 U173 ( .B1(n90), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U174 ( .B1(n90), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X2 U175 ( .B1(n46), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X2 U176 ( .B1(n46), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U177 ( .B1(n71), .B2(n84), .A(n72), .ZN(n70) );
  OAI21_X2 U178 ( .B1(n73), .B2(n79), .A(n74), .ZN(n72) );
  AOI21_X2 U179 ( .B1(n211), .B2(n43), .A(n38), .ZN(n36) );
  AOI21_X2 U180 ( .B1(n113), .B2(n121), .A(n114), .ZN(n112) );
  NOR2_X2 U181 ( .A1(n118), .A2(n115), .ZN(n113) );
  OAI21_X2 U182 ( .B1(n115), .B2(n119), .A(n116), .ZN(n114) );
  OAI21_X2 U183 ( .B1(n36), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X2 U184 ( .B1(n62), .B2(n66), .A(n63), .ZN(n61) );
  OAI21_X2 U185 ( .B1(n104), .B2(n110), .A(n105), .ZN(n103) );
  OAI21_X2 U186 ( .B1(n112), .B2(n92), .A(n93), .ZN(n91) );
  AOI21_X2 U187 ( .B1(n94), .B2(n103), .A(n95), .ZN(n93) );
  NOR2_X2 U188 ( .A1(n99), .A2(n96), .ZN(n94) );
  AOI21_X2 U189 ( .B1(n52), .B2(n61), .A(n53), .ZN(n51) );
  OAI21_X2 U190 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  AOI21_X2 U191 ( .B1(n29), .B2(n213), .A(n24), .ZN(n22) );
  AOI21_X2 U192 ( .B1(n80), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X2 U193 ( .B1(n46), .B2(n212), .A(n43), .ZN(n41) );
  OAI21_X2 U194 ( .B1(n122), .B2(n124), .A(n123), .ZN(n121) );
  OAI21_X2 U195 ( .B1(n85), .B2(n89), .A(n86), .ZN(n84) );
  OAI21_X2 U196 ( .B1(n96), .B2(n100), .A(n97), .ZN(n95) );
  OAI21_X2 U197 ( .B1(n101), .B2(n99), .A(n100), .ZN(n98) );
  OAI21_X2 U198 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X2 U199 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NOR2_X2 U200 ( .A1(n57), .A2(n54), .ZN(n52) );
  NOR2_X2 U201 ( .A1(n78), .A2(n73), .ZN(n71) );
  NOR2_X2 U202 ( .A1(n109), .A2(n104), .ZN(n102) );
  NOR2_X2 U203 ( .A1(n65), .A2(n62), .ZN(n60) );
  NOR2_X2 U204 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U205 ( .A1(n88), .A2(n85), .ZN(n83) );
  AOI21_X2 U206 ( .B1(n111), .B2(n140), .A(n108), .ZN(n106) );
  OAI21_X2 U207 ( .B1(n120), .B2(n118), .A(n119), .ZN(n117) );
  OAI21_X2 U208 ( .B1(n90), .B2(n88), .A(n89), .ZN(n87) );
  NOR2_X2 U209 ( .A1(A[3]), .A2(B[3]), .ZN(n115) );
  NOR2_X2 U210 ( .A1(A[7]), .A2(B[7]), .ZN(n96) );
  NOR2_X2 U211 ( .A1(A[5]), .A2(B[5]), .ZN(n104) );
  NOR2_X2 U212 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  NOR2_X2 U213 ( .A1(A[13]), .A2(B[13]), .ZN(n62) );
  NOR2_X2 U214 ( .A1(A[11]), .A2(B[11]), .ZN(n73) );
  NOR2_X2 U215 ( .A1(A[9]), .A2(B[9]), .ZN(n85) );
  NOR2_X2 U216 ( .A1(A[18]), .A2(B[18]), .ZN(n30) );
  NOR2_X2 U217 ( .A1(A[2]), .A2(B[2]), .ZN(n118) );
  NOR2_X2 U218 ( .A1(A[6]), .A2(B[6]), .ZN(n99) );
  NOR2_X2 U219 ( .A1(A[8]), .A2(B[8]), .ZN(n88) );
  NOR2_X2 U220 ( .A1(A[12]), .A2(B[12]), .ZN(n65) );
  NOR2_X2 U221 ( .A1(A[14]), .A2(B[14]), .ZN(n57) );
  NOR2_X2 U222 ( .A1(A[1]), .A2(B[1]), .ZN(n122) );
  NOR2_X2 U223 ( .A1(A[0]), .A2(B[0]), .ZN(n124) );
  NOR2_X2 U224 ( .A1(A[4]), .A2(B[4]), .ZN(n109) );
  NOR2_X2 U225 ( .A1(A[10]), .A2(B[10]), .ZN(n78) );
  OAI21_X2 U226 ( .B1(n47), .B2(n21), .A(n22), .ZN(CO) );
  OR2_X1 U227 ( .A1(A[17]), .A2(B[17]), .ZN(n211) );
  OR2_X1 U228 ( .A1(A[16]), .A2(B[16]), .ZN(n212) );
  OR2_X1 U229 ( .A1(A[19]), .A2(B[19]), .ZN(n213) );
  INV_X4 U230 ( .A(n91), .ZN(n90) );
  INV_X4 U231 ( .A(n84), .ZN(n82) );
  INV_X4 U232 ( .A(n83), .ZN(n81) );
  INV_X4 U233 ( .A(n79), .ZN(n77) );
  INV_X4 U234 ( .A(n68), .ZN(n67) );
  INV_X4 U235 ( .A(n47), .ZN(n46) );
  INV_X4 U236 ( .A(n45), .ZN(n43) );
  INV_X4 U237 ( .A(n40), .ZN(n38) );
  INV_X4 U238 ( .A(n36), .ZN(n34) );
  INV_X4 U239 ( .A(n35), .ZN(n33) );
  INV_X4 U240 ( .A(n26), .ZN(n24) );
  INV_X4 U241 ( .A(n122), .ZN(n143) );
  INV_X4 U242 ( .A(n118), .ZN(n142) );
  INV_X4 U243 ( .A(n115), .ZN(n141) );
  INV_X4 U244 ( .A(n104), .ZN(n139) );
  INV_X4 U245 ( .A(n99), .ZN(n138) );
  INV_X4 U246 ( .A(n96), .ZN(n137) );
  INV_X4 U247 ( .A(n88), .ZN(n136) );
  INV_X4 U248 ( .A(n85), .ZN(n135) );
  INV_X4 U249 ( .A(n78), .ZN(n76) );
  INV_X4 U250 ( .A(n73), .ZN(n133) );
  INV_X4 U251 ( .A(n65), .ZN(n132) );
  INV_X4 U252 ( .A(n62), .ZN(n131) );
  INV_X4 U253 ( .A(n57), .ZN(n130) );
  INV_X4 U254 ( .A(n54), .ZN(n129) );
  INV_X4 U255 ( .A(n30), .ZN(n126) );
  INV_X4 U256 ( .A(n121), .ZN(n120) );
  INV_X4 U257 ( .A(n112), .ZN(n111) );
  INV_X4 U258 ( .A(n110), .ZN(n108) );
  INV_X4 U259 ( .A(n109), .ZN(n140) );
endmodule


module pipleline_stage_5 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n105;
  wire   [20:0] stage_result;

  pipleline_stage_5_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(stage_out[0]) );
  INV_X4 U6 ( .A(n105), .ZN(q) );
  BUF_X4 U7 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U8 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U9 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U10 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U11 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U12 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U13 ( .A(divided[0]), .Z(stage_out[1]) );
  XNOR2_X2 U14 ( .A(divided[27]), .B(stage_result[20]), .ZN(n105) );
  MUX2_X2 U15 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U16 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U17 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U18 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U19 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U20 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U22 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U23 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U24 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U25 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U26 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U27 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U28 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U29 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U30 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U31 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U32 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U33 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U34 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n38, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n129, n130, n131,
         n132, n133, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n211, n212, n213;

  XOR2_X2 U2 ( .A(n1), .B(n27), .Z(SUM[19]) );
  NAND2_X2 U4 ( .A1(n28), .A2(n213), .ZN(n21) );
  NAND2_X2 U8 ( .A1(n213), .A2(n26), .ZN(n1) );
  NAND2_X2 U11 ( .A1(A[19]), .A2(B[19]), .ZN(n26) );
  XOR2_X2 U12 ( .A(n2), .B(n32), .Z(SUM[18]) );
  NAND2_X2 U16 ( .A1(n126), .A2(n31), .ZN(n2) );
  NAND2_X2 U19 ( .A1(A[18]), .A2(B[18]), .ZN(n31) );
  XOR2_X2 U20 ( .A(n3), .B(n41), .Z(SUM[17]) );
  NAND2_X2 U24 ( .A1(n212), .A2(n211), .ZN(n35) );
  NAND2_X2 U28 ( .A1(n211), .A2(n40), .ZN(n3) );
  NAND2_X2 U31 ( .A1(A[17]), .A2(B[17]), .ZN(n40) );
  XNOR2_X2 U32 ( .A(n46), .B(n4), .ZN(SUM[16]) );
  NAND2_X2 U36 ( .A1(n212), .A2(n45), .ZN(n4) );
  NAND2_X2 U39 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U40 ( .A(n56), .B(n5), .ZN(SUM[15]) );
  NAND2_X2 U45 ( .A1(n60), .A2(n52), .ZN(n50) );
  NAND2_X2 U49 ( .A1(n129), .A2(n55), .ZN(n5) );
  NAND2_X2 U52 ( .A1(A[15]), .A2(B[15]), .ZN(n55) );
  XOR2_X2 U53 ( .A(n6), .B(n59), .Z(SUM[14]) );
  NAND2_X2 U55 ( .A1(n130), .A2(n58), .ZN(n6) );
  NAND2_X2 U58 ( .A1(A[14]), .A2(B[14]), .ZN(n58) );
  XNOR2_X2 U59 ( .A(n64), .B(n7), .ZN(SUM[13]) );
  NAND2_X2 U63 ( .A1(n131), .A2(n63), .ZN(n7) );
  NAND2_X2 U66 ( .A1(A[13]), .A2(B[13]), .ZN(n63) );
  XOR2_X2 U67 ( .A(n8), .B(n67), .Z(SUM[12]) );
  NAND2_X2 U69 ( .A1(n132), .A2(n66), .ZN(n8) );
  NAND2_X2 U72 ( .A1(A[12]), .A2(B[12]), .ZN(n66) );
  XOR2_X2 U73 ( .A(n9), .B(n75), .Z(SUM[11]) );
  NAND2_X2 U76 ( .A1(n83), .A2(n71), .ZN(n69) );
  NAND2_X2 U80 ( .A1(n133), .A2(n74), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[11]), .A2(B[11]), .ZN(n74) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[10]) );
  NAND2_X2 U88 ( .A1(n76), .A2(n79), .ZN(n10) );
  NAND2_X2 U91 ( .A1(A[10]), .A2(B[10]), .ZN(n79) );
  XNOR2_X2 U92 ( .A(n87), .B(n11), .ZN(SUM[9]) );
  NAND2_X2 U98 ( .A1(n135), .A2(n86), .ZN(n11) );
  NAND2_X2 U101 ( .A1(A[9]), .A2(B[9]), .ZN(n86) );
  XOR2_X2 U102 ( .A(n12), .B(n90), .Z(SUM[8]) );
  NAND2_X2 U104 ( .A1(n136), .A2(n89), .ZN(n12) );
  NAND2_X2 U107 ( .A1(A[8]), .A2(B[8]), .ZN(n89) );
  XNOR2_X2 U108 ( .A(n98), .B(n13), .ZN(SUM[7]) );
  NAND2_X2 U111 ( .A1(n102), .A2(n94), .ZN(n92) );
  NAND2_X2 U115 ( .A1(n137), .A2(n97), .ZN(n13) );
  NAND2_X2 U118 ( .A1(A[7]), .A2(B[7]), .ZN(n97) );
  XOR2_X2 U119 ( .A(n14), .B(n101), .Z(SUM[6]) );
  NAND2_X2 U121 ( .A1(n138), .A2(n100), .ZN(n14) );
  NAND2_X2 U124 ( .A1(A[6]), .A2(B[6]), .ZN(n100) );
  XOR2_X2 U125 ( .A(n15), .B(n106), .Z(SUM[5]) );
  NAND2_X2 U129 ( .A1(n139), .A2(n105), .ZN(n15) );
  NAND2_X2 U132 ( .A1(A[5]), .A2(B[5]), .ZN(n105) );
  XNOR2_X2 U133 ( .A(n111), .B(n16), .ZN(SUM[4]) );
  NAND2_X2 U137 ( .A1(n140), .A2(n110), .ZN(n16) );
  NAND2_X2 U140 ( .A1(A[4]), .A2(B[4]), .ZN(n110) );
  XNOR2_X2 U141 ( .A(n117), .B(n17), .ZN(SUM[3]) );
  NAND2_X2 U146 ( .A1(n141), .A2(n116), .ZN(n17) );
  NAND2_X2 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n116) );
  XOR2_X2 U150 ( .A(n18), .B(n120), .Z(SUM[2]) );
  NAND2_X2 U152 ( .A1(n142), .A2(n119), .ZN(n18) );
  NAND2_X2 U155 ( .A1(A[2]), .A2(B[2]), .ZN(n119) );
  XOR2_X2 U156 ( .A(n124), .B(n19), .Z(SUM[1]) );
  NAND2_X2 U159 ( .A1(n143), .A2(n123), .ZN(n19) );
  NAND2_X2 U162 ( .A1(A[1]), .A2(B[1]), .ZN(n123) );
  XNOR2_X2 U163 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U168 ( .B1(n111), .B2(n102), .A(n103), .ZN(n101) );
  AOI21_X2 U169 ( .B1(n68), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X2 U170 ( .B1(n91), .B2(n48), .A(n49), .ZN(n47) );
  NOR2_X2 U171 ( .A1(n69), .A2(n50), .ZN(n48) );
  OAI21_X2 U172 ( .B1(n70), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X2 U173 ( .B1(n90), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U174 ( .B1(n90), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X2 U175 ( .B1(n46), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X2 U176 ( .B1(n46), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U177 ( .B1(n71), .B2(n84), .A(n72), .ZN(n70) );
  OAI21_X2 U178 ( .B1(n73), .B2(n79), .A(n74), .ZN(n72) );
  AOI21_X2 U179 ( .B1(n211), .B2(n43), .A(n38), .ZN(n36) );
  AOI21_X2 U180 ( .B1(n113), .B2(n121), .A(n114), .ZN(n112) );
  NOR2_X2 U181 ( .A1(n118), .A2(n115), .ZN(n113) );
  OAI21_X2 U182 ( .B1(n115), .B2(n119), .A(n116), .ZN(n114) );
  OAI21_X2 U183 ( .B1(n36), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X2 U184 ( .B1(n62), .B2(n66), .A(n63), .ZN(n61) );
  OAI21_X2 U185 ( .B1(n104), .B2(n110), .A(n105), .ZN(n103) );
  OAI21_X2 U186 ( .B1(n112), .B2(n92), .A(n93), .ZN(n91) );
  AOI21_X2 U187 ( .B1(n94), .B2(n103), .A(n95), .ZN(n93) );
  NOR2_X2 U188 ( .A1(n99), .A2(n96), .ZN(n94) );
  AOI21_X2 U189 ( .B1(n52), .B2(n61), .A(n53), .ZN(n51) );
  OAI21_X2 U190 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  AOI21_X2 U191 ( .B1(n29), .B2(n213), .A(n24), .ZN(n22) );
  AOI21_X2 U192 ( .B1(n80), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X2 U193 ( .B1(n46), .B2(n212), .A(n43), .ZN(n41) );
  OAI21_X2 U194 ( .B1(n122), .B2(n124), .A(n123), .ZN(n121) );
  OAI21_X2 U195 ( .B1(n85), .B2(n89), .A(n86), .ZN(n84) );
  OAI21_X2 U196 ( .B1(n96), .B2(n100), .A(n97), .ZN(n95) );
  OAI21_X2 U197 ( .B1(n101), .B2(n99), .A(n100), .ZN(n98) );
  OAI21_X2 U198 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X2 U199 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NOR2_X2 U200 ( .A1(n57), .A2(n54), .ZN(n52) );
  NOR2_X2 U201 ( .A1(n78), .A2(n73), .ZN(n71) );
  NOR2_X2 U202 ( .A1(n109), .A2(n104), .ZN(n102) );
  NOR2_X2 U203 ( .A1(n65), .A2(n62), .ZN(n60) );
  NOR2_X2 U204 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U205 ( .A1(n88), .A2(n85), .ZN(n83) );
  AOI21_X2 U206 ( .B1(n111), .B2(n140), .A(n108), .ZN(n106) );
  OAI21_X2 U207 ( .B1(n120), .B2(n118), .A(n119), .ZN(n117) );
  OAI21_X2 U208 ( .B1(n90), .B2(n88), .A(n89), .ZN(n87) );
  NOR2_X2 U209 ( .A1(A[3]), .A2(B[3]), .ZN(n115) );
  NOR2_X2 U210 ( .A1(A[7]), .A2(B[7]), .ZN(n96) );
  NOR2_X2 U211 ( .A1(A[5]), .A2(B[5]), .ZN(n104) );
  NOR2_X2 U212 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  NOR2_X2 U213 ( .A1(A[13]), .A2(B[13]), .ZN(n62) );
  NOR2_X2 U214 ( .A1(A[11]), .A2(B[11]), .ZN(n73) );
  NOR2_X2 U215 ( .A1(A[9]), .A2(B[9]), .ZN(n85) );
  NOR2_X2 U216 ( .A1(A[18]), .A2(B[18]), .ZN(n30) );
  NOR2_X2 U217 ( .A1(A[2]), .A2(B[2]), .ZN(n118) );
  NOR2_X2 U218 ( .A1(A[6]), .A2(B[6]), .ZN(n99) );
  NOR2_X2 U219 ( .A1(A[8]), .A2(B[8]), .ZN(n88) );
  NOR2_X2 U220 ( .A1(A[12]), .A2(B[12]), .ZN(n65) );
  NOR2_X2 U221 ( .A1(A[14]), .A2(B[14]), .ZN(n57) );
  NOR2_X2 U222 ( .A1(A[1]), .A2(B[1]), .ZN(n122) );
  NOR2_X2 U223 ( .A1(A[0]), .A2(B[0]), .ZN(n124) );
  NOR2_X2 U224 ( .A1(A[4]), .A2(B[4]), .ZN(n109) );
  NOR2_X2 U225 ( .A1(A[10]), .A2(B[10]), .ZN(n78) );
  OAI21_X2 U226 ( .B1(n47), .B2(n21), .A(n22), .ZN(CO) );
  OR2_X1 U227 ( .A1(A[17]), .A2(B[17]), .ZN(n211) );
  OR2_X1 U228 ( .A1(A[16]), .A2(B[16]), .ZN(n212) );
  OR2_X1 U229 ( .A1(A[19]), .A2(B[19]), .ZN(n213) );
  INV_X4 U230 ( .A(n91), .ZN(n90) );
  INV_X4 U231 ( .A(n84), .ZN(n82) );
  INV_X4 U232 ( .A(n83), .ZN(n81) );
  INV_X4 U233 ( .A(n79), .ZN(n77) );
  INV_X4 U234 ( .A(n68), .ZN(n67) );
  INV_X4 U235 ( .A(n47), .ZN(n46) );
  INV_X4 U236 ( .A(n45), .ZN(n43) );
  INV_X4 U237 ( .A(n40), .ZN(n38) );
  INV_X4 U238 ( .A(n36), .ZN(n34) );
  INV_X4 U239 ( .A(n35), .ZN(n33) );
  INV_X4 U240 ( .A(n26), .ZN(n24) );
  INV_X4 U241 ( .A(n122), .ZN(n143) );
  INV_X4 U242 ( .A(n118), .ZN(n142) );
  INV_X4 U243 ( .A(n115), .ZN(n141) );
  INV_X4 U244 ( .A(n104), .ZN(n139) );
  INV_X4 U245 ( .A(n99), .ZN(n138) );
  INV_X4 U246 ( .A(n96), .ZN(n137) );
  INV_X4 U247 ( .A(n88), .ZN(n136) );
  INV_X4 U248 ( .A(n85), .ZN(n135) );
  INV_X4 U249 ( .A(n78), .ZN(n76) );
  INV_X4 U250 ( .A(n73), .ZN(n133) );
  INV_X4 U251 ( .A(n65), .ZN(n132) );
  INV_X4 U252 ( .A(n62), .ZN(n131) );
  INV_X4 U253 ( .A(n57), .ZN(n130) );
  INV_X4 U254 ( .A(n54), .ZN(n129) );
  INV_X4 U255 ( .A(n30), .ZN(n126) );
  INV_X4 U256 ( .A(n121), .ZN(n120) );
  INV_X4 U257 ( .A(n112), .ZN(n111) );
  INV_X4 U258 ( .A(n110), .ZN(n108) );
  INV_X4 U259 ( .A(n109), .ZN(n140) );
endmodule


module pipleline_stage_4 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n105;
  wire   [20:0] stage_result;

  pipleline_stage_4_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(stage_out[0]) );
  INV_X4 U6 ( .A(n105), .ZN(q) );
  BUF_X4 U7 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U8 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U9 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U10 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U11 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U12 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U13 ( .A(divided[0]), .Z(stage_out[1]) );
  XNOR2_X2 U14 ( .A(divided[27]), .B(stage_result[20]), .ZN(n105) );
  MUX2_X2 U15 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U16 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U17 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U18 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U19 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U20 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U22 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U23 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U24 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U25 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U26 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U27 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U28 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U29 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U30 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U31 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U32 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U33 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U34 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n38, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n129, n130, n131,
         n132, n133, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n211, n212, n213;

  XOR2_X2 U2 ( .A(n1), .B(n27), .Z(SUM[19]) );
  NAND2_X2 U4 ( .A1(n28), .A2(n213), .ZN(n21) );
  NAND2_X2 U8 ( .A1(n213), .A2(n26), .ZN(n1) );
  NAND2_X2 U11 ( .A1(A[19]), .A2(B[19]), .ZN(n26) );
  XOR2_X2 U12 ( .A(n2), .B(n32), .Z(SUM[18]) );
  NAND2_X2 U16 ( .A1(n126), .A2(n31), .ZN(n2) );
  NAND2_X2 U19 ( .A1(A[18]), .A2(B[18]), .ZN(n31) );
  XOR2_X2 U20 ( .A(n3), .B(n41), .Z(SUM[17]) );
  NAND2_X2 U24 ( .A1(n212), .A2(n211), .ZN(n35) );
  NAND2_X2 U28 ( .A1(n211), .A2(n40), .ZN(n3) );
  NAND2_X2 U31 ( .A1(A[17]), .A2(B[17]), .ZN(n40) );
  XNOR2_X2 U32 ( .A(n46), .B(n4), .ZN(SUM[16]) );
  NAND2_X2 U36 ( .A1(n212), .A2(n45), .ZN(n4) );
  NAND2_X2 U39 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U40 ( .A(n56), .B(n5), .ZN(SUM[15]) );
  NAND2_X2 U45 ( .A1(n60), .A2(n52), .ZN(n50) );
  NAND2_X2 U49 ( .A1(n129), .A2(n55), .ZN(n5) );
  NAND2_X2 U52 ( .A1(A[15]), .A2(B[15]), .ZN(n55) );
  XOR2_X2 U53 ( .A(n6), .B(n59), .Z(SUM[14]) );
  NAND2_X2 U55 ( .A1(n130), .A2(n58), .ZN(n6) );
  NAND2_X2 U58 ( .A1(A[14]), .A2(B[14]), .ZN(n58) );
  XNOR2_X2 U59 ( .A(n64), .B(n7), .ZN(SUM[13]) );
  NAND2_X2 U63 ( .A1(n131), .A2(n63), .ZN(n7) );
  NAND2_X2 U66 ( .A1(A[13]), .A2(B[13]), .ZN(n63) );
  XOR2_X2 U67 ( .A(n8), .B(n67), .Z(SUM[12]) );
  NAND2_X2 U69 ( .A1(n132), .A2(n66), .ZN(n8) );
  NAND2_X2 U72 ( .A1(A[12]), .A2(B[12]), .ZN(n66) );
  XOR2_X2 U73 ( .A(n9), .B(n75), .Z(SUM[11]) );
  NAND2_X2 U76 ( .A1(n83), .A2(n71), .ZN(n69) );
  NAND2_X2 U80 ( .A1(n133), .A2(n74), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[11]), .A2(B[11]), .ZN(n74) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[10]) );
  NAND2_X2 U88 ( .A1(n76), .A2(n79), .ZN(n10) );
  NAND2_X2 U91 ( .A1(A[10]), .A2(B[10]), .ZN(n79) );
  XNOR2_X2 U92 ( .A(n87), .B(n11), .ZN(SUM[9]) );
  NAND2_X2 U98 ( .A1(n135), .A2(n86), .ZN(n11) );
  NAND2_X2 U101 ( .A1(A[9]), .A2(B[9]), .ZN(n86) );
  XOR2_X2 U102 ( .A(n12), .B(n90), .Z(SUM[8]) );
  NAND2_X2 U104 ( .A1(n136), .A2(n89), .ZN(n12) );
  NAND2_X2 U107 ( .A1(A[8]), .A2(B[8]), .ZN(n89) );
  XNOR2_X2 U108 ( .A(n98), .B(n13), .ZN(SUM[7]) );
  NAND2_X2 U111 ( .A1(n102), .A2(n94), .ZN(n92) );
  NAND2_X2 U115 ( .A1(n137), .A2(n97), .ZN(n13) );
  NAND2_X2 U118 ( .A1(A[7]), .A2(B[7]), .ZN(n97) );
  XOR2_X2 U119 ( .A(n14), .B(n101), .Z(SUM[6]) );
  NAND2_X2 U121 ( .A1(n138), .A2(n100), .ZN(n14) );
  NAND2_X2 U124 ( .A1(A[6]), .A2(B[6]), .ZN(n100) );
  XOR2_X2 U125 ( .A(n15), .B(n106), .Z(SUM[5]) );
  NAND2_X2 U129 ( .A1(n139), .A2(n105), .ZN(n15) );
  NAND2_X2 U132 ( .A1(A[5]), .A2(B[5]), .ZN(n105) );
  XNOR2_X2 U133 ( .A(n111), .B(n16), .ZN(SUM[4]) );
  NAND2_X2 U137 ( .A1(n140), .A2(n110), .ZN(n16) );
  NAND2_X2 U140 ( .A1(A[4]), .A2(B[4]), .ZN(n110) );
  XNOR2_X2 U141 ( .A(n117), .B(n17), .ZN(SUM[3]) );
  NAND2_X2 U146 ( .A1(n141), .A2(n116), .ZN(n17) );
  NAND2_X2 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n116) );
  XOR2_X2 U150 ( .A(n18), .B(n120), .Z(SUM[2]) );
  NAND2_X2 U152 ( .A1(n142), .A2(n119), .ZN(n18) );
  NAND2_X2 U155 ( .A1(A[2]), .A2(B[2]), .ZN(n119) );
  XOR2_X2 U156 ( .A(n124), .B(n19), .Z(SUM[1]) );
  NAND2_X2 U159 ( .A1(n143), .A2(n123), .ZN(n19) );
  NAND2_X2 U162 ( .A1(A[1]), .A2(B[1]), .ZN(n123) );
  XNOR2_X2 U163 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U168 ( .B1(n111), .B2(n102), .A(n103), .ZN(n101) );
  AOI21_X2 U169 ( .B1(n68), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X2 U170 ( .B1(n91), .B2(n48), .A(n49), .ZN(n47) );
  NOR2_X2 U171 ( .A1(n69), .A2(n50), .ZN(n48) );
  OAI21_X2 U172 ( .B1(n70), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X2 U173 ( .B1(n90), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U174 ( .B1(n90), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X2 U175 ( .B1(n46), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X2 U176 ( .B1(n46), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U177 ( .B1(n71), .B2(n84), .A(n72), .ZN(n70) );
  OAI21_X2 U178 ( .B1(n73), .B2(n79), .A(n74), .ZN(n72) );
  AOI21_X2 U179 ( .B1(n211), .B2(n43), .A(n38), .ZN(n36) );
  AOI21_X2 U180 ( .B1(n113), .B2(n121), .A(n114), .ZN(n112) );
  NOR2_X2 U181 ( .A1(n118), .A2(n115), .ZN(n113) );
  OAI21_X2 U182 ( .B1(n115), .B2(n119), .A(n116), .ZN(n114) );
  OAI21_X2 U183 ( .B1(n36), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X2 U184 ( .B1(n62), .B2(n66), .A(n63), .ZN(n61) );
  OAI21_X2 U185 ( .B1(n104), .B2(n110), .A(n105), .ZN(n103) );
  OAI21_X2 U186 ( .B1(n112), .B2(n92), .A(n93), .ZN(n91) );
  AOI21_X2 U187 ( .B1(n94), .B2(n103), .A(n95), .ZN(n93) );
  NOR2_X2 U188 ( .A1(n99), .A2(n96), .ZN(n94) );
  AOI21_X2 U189 ( .B1(n52), .B2(n61), .A(n53), .ZN(n51) );
  OAI21_X2 U190 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  AOI21_X2 U191 ( .B1(n29), .B2(n213), .A(n24), .ZN(n22) );
  AOI21_X2 U192 ( .B1(n80), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X2 U193 ( .B1(n46), .B2(n212), .A(n43), .ZN(n41) );
  OAI21_X2 U194 ( .B1(n122), .B2(n124), .A(n123), .ZN(n121) );
  OAI21_X2 U195 ( .B1(n85), .B2(n89), .A(n86), .ZN(n84) );
  OAI21_X2 U196 ( .B1(n96), .B2(n100), .A(n97), .ZN(n95) );
  OAI21_X2 U197 ( .B1(n101), .B2(n99), .A(n100), .ZN(n98) );
  OAI21_X2 U198 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X2 U199 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NOR2_X2 U200 ( .A1(n57), .A2(n54), .ZN(n52) );
  NOR2_X2 U201 ( .A1(n78), .A2(n73), .ZN(n71) );
  NOR2_X2 U202 ( .A1(n109), .A2(n104), .ZN(n102) );
  NOR2_X2 U203 ( .A1(n65), .A2(n62), .ZN(n60) );
  NOR2_X2 U204 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U205 ( .A1(n88), .A2(n85), .ZN(n83) );
  AOI21_X2 U206 ( .B1(n111), .B2(n140), .A(n108), .ZN(n106) );
  OAI21_X2 U207 ( .B1(n120), .B2(n118), .A(n119), .ZN(n117) );
  OAI21_X2 U208 ( .B1(n90), .B2(n88), .A(n89), .ZN(n87) );
  NOR2_X2 U209 ( .A1(A[3]), .A2(B[3]), .ZN(n115) );
  NOR2_X2 U210 ( .A1(A[7]), .A2(B[7]), .ZN(n96) );
  NOR2_X2 U211 ( .A1(A[5]), .A2(B[5]), .ZN(n104) );
  NOR2_X2 U212 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  NOR2_X2 U213 ( .A1(A[13]), .A2(B[13]), .ZN(n62) );
  NOR2_X2 U214 ( .A1(A[11]), .A2(B[11]), .ZN(n73) );
  NOR2_X2 U215 ( .A1(A[9]), .A2(B[9]), .ZN(n85) );
  NOR2_X2 U216 ( .A1(A[18]), .A2(B[18]), .ZN(n30) );
  NOR2_X2 U217 ( .A1(A[2]), .A2(B[2]), .ZN(n118) );
  NOR2_X2 U218 ( .A1(A[6]), .A2(B[6]), .ZN(n99) );
  NOR2_X2 U219 ( .A1(A[8]), .A2(B[8]), .ZN(n88) );
  NOR2_X2 U220 ( .A1(A[12]), .A2(B[12]), .ZN(n65) );
  NOR2_X2 U221 ( .A1(A[14]), .A2(B[14]), .ZN(n57) );
  NOR2_X2 U222 ( .A1(A[1]), .A2(B[1]), .ZN(n122) );
  NOR2_X2 U223 ( .A1(A[0]), .A2(B[0]), .ZN(n124) );
  NOR2_X2 U224 ( .A1(A[4]), .A2(B[4]), .ZN(n109) );
  NOR2_X2 U225 ( .A1(A[10]), .A2(B[10]), .ZN(n78) );
  OAI21_X2 U226 ( .B1(n47), .B2(n21), .A(n22), .ZN(CO) );
  OR2_X1 U227 ( .A1(A[17]), .A2(B[17]), .ZN(n211) );
  OR2_X1 U228 ( .A1(A[16]), .A2(B[16]), .ZN(n212) );
  OR2_X1 U229 ( .A1(A[19]), .A2(B[19]), .ZN(n213) );
  INV_X4 U230 ( .A(n91), .ZN(n90) );
  INV_X4 U231 ( .A(n84), .ZN(n82) );
  INV_X4 U232 ( .A(n83), .ZN(n81) );
  INV_X4 U233 ( .A(n79), .ZN(n77) );
  INV_X4 U234 ( .A(n68), .ZN(n67) );
  INV_X4 U235 ( .A(n47), .ZN(n46) );
  INV_X4 U236 ( .A(n45), .ZN(n43) );
  INV_X4 U237 ( .A(n40), .ZN(n38) );
  INV_X4 U238 ( .A(n36), .ZN(n34) );
  INV_X4 U239 ( .A(n35), .ZN(n33) );
  INV_X4 U240 ( .A(n26), .ZN(n24) );
  INV_X4 U241 ( .A(n122), .ZN(n143) );
  INV_X4 U242 ( .A(n118), .ZN(n142) );
  INV_X4 U243 ( .A(n115), .ZN(n141) );
  INV_X4 U244 ( .A(n104), .ZN(n139) );
  INV_X4 U245 ( .A(n99), .ZN(n138) );
  INV_X4 U246 ( .A(n96), .ZN(n137) );
  INV_X4 U247 ( .A(n88), .ZN(n136) );
  INV_X4 U248 ( .A(n85), .ZN(n135) );
  INV_X4 U249 ( .A(n78), .ZN(n76) );
  INV_X4 U250 ( .A(n73), .ZN(n133) );
  INV_X4 U251 ( .A(n65), .ZN(n132) );
  INV_X4 U252 ( .A(n62), .ZN(n131) );
  INV_X4 U253 ( .A(n57), .ZN(n130) );
  INV_X4 U254 ( .A(n54), .ZN(n129) );
  INV_X4 U255 ( .A(n30), .ZN(n126) );
  INV_X4 U256 ( .A(n121), .ZN(n120) );
  INV_X4 U257 ( .A(n112), .ZN(n111) );
  INV_X4 U258 ( .A(n110), .ZN(n108) );
  INV_X4 U259 ( .A(n109), .ZN(n140) );
endmodule


module pipleline_stage_3 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n105;
  wire   [20:0] stage_result;

  pipleline_stage_3_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(stage_out[0]) );
  INV_X4 U6 ( .A(n105), .ZN(q) );
  BUF_X4 U7 ( .A(divided[0]), .Z(stage_out[1]) );
  BUF_X4 U8 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U9 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U10 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U11 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U12 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U13 ( .A(divided[6]), .Z(stage_out[7]) );
  XNOR2_X2 U14 ( .A(divided[27]), .B(stage_result[20]), .ZN(n105) );
  MUX2_X2 U15 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U16 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U17 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U18 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U19 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U20 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U22 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U23 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U24 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U25 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U26 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U27 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U28 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U29 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U30 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U31 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U32 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U33 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U34 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n24, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n38, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n129, n130, n131,
         n132, n133, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n211, n212, n213;

  XOR2_X2 U2 ( .A(n1), .B(n27), .Z(SUM[19]) );
  NAND2_X2 U4 ( .A1(n28), .A2(n213), .ZN(n21) );
  NAND2_X2 U8 ( .A1(n213), .A2(n26), .ZN(n1) );
  NAND2_X2 U11 ( .A1(A[19]), .A2(B[19]), .ZN(n26) );
  XOR2_X2 U12 ( .A(n2), .B(n32), .Z(SUM[18]) );
  NAND2_X2 U16 ( .A1(n126), .A2(n31), .ZN(n2) );
  NAND2_X2 U19 ( .A1(A[18]), .A2(B[18]), .ZN(n31) );
  XOR2_X2 U20 ( .A(n3), .B(n41), .Z(SUM[17]) );
  NAND2_X2 U24 ( .A1(n212), .A2(n211), .ZN(n35) );
  NAND2_X2 U28 ( .A1(n211), .A2(n40), .ZN(n3) );
  NAND2_X2 U31 ( .A1(A[17]), .A2(B[17]), .ZN(n40) );
  XNOR2_X2 U32 ( .A(n46), .B(n4), .ZN(SUM[16]) );
  NAND2_X2 U36 ( .A1(n212), .A2(n45), .ZN(n4) );
  NAND2_X2 U39 ( .A1(A[16]), .A2(B[16]), .ZN(n45) );
  XNOR2_X2 U40 ( .A(n56), .B(n5), .ZN(SUM[15]) );
  NAND2_X2 U45 ( .A1(n60), .A2(n52), .ZN(n50) );
  NAND2_X2 U49 ( .A1(n129), .A2(n55), .ZN(n5) );
  NAND2_X2 U52 ( .A1(A[15]), .A2(B[15]), .ZN(n55) );
  XOR2_X2 U53 ( .A(n6), .B(n59), .Z(SUM[14]) );
  NAND2_X2 U55 ( .A1(n130), .A2(n58), .ZN(n6) );
  NAND2_X2 U58 ( .A1(A[14]), .A2(B[14]), .ZN(n58) );
  XNOR2_X2 U59 ( .A(n64), .B(n7), .ZN(SUM[13]) );
  NAND2_X2 U63 ( .A1(n131), .A2(n63), .ZN(n7) );
  NAND2_X2 U66 ( .A1(A[13]), .A2(B[13]), .ZN(n63) );
  XOR2_X2 U67 ( .A(n8), .B(n67), .Z(SUM[12]) );
  NAND2_X2 U69 ( .A1(n132), .A2(n66), .ZN(n8) );
  NAND2_X2 U72 ( .A1(A[12]), .A2(B[12]), .ZN(n66) );
  XOR2_X2 U73 ( .A(n9), .B(n75), .Z(SUM[11]) );
  NAND2_X2 U76 ( .A1(n83), .A2(n71), .ZN(n69) );
  NAND2_X2 U80 ( .A1(n133), .A2(n74), .ZN(n9) );
  NAND2_X2 U83 ( .A1(A[11]), .A2(B[11]), .ZN(n74) );
  XNOR2_X2 U84 ( .A(n80), .B(n10), .ZN(SUM[10]) );
  NAND2_X2 U88 ( .A1(n76), .A2(n79), .ZN(n10) );
  NAND2_X2 U91 ( .A1(A[10]), .A2(B[10]), .ZN(n79) );
  XNOR2_X2 U92 ( .A(n87), .B(n11), .ZN(SUM[9]) );
  NAND2_X2 U98 ( .A1(n135), .A2(n86), .ZN(n11) );
  NAND2_X2 U101 ( .A1(A[9]), .A2(B[9]), .ZN(n86) );
  XOR2_X2 U102 ( .A(n12), .B(n90), .Z(SUM[8]) );
  NAND2_X2 U104 ( .A1(n136), .A2(n89), .ZN(n12) );
  NAND2_X2 U107 ( .A1(A[8]), .A2(B[8]), .ZN(n89) );
  XNOR2_X2 U108 ( .A(n98), .B(n13), .ZN(SUM[7]) );
  NAND2_X2 U111 ( .A1(n102), .A2(n94), .ZN(n92) );
  NAND2_X2 U115 ( .A1(n137), .A2(n97), .ZN(n13) );
  NAND2_X2 U118 ( .A1(A[7]), .A2(B[7]), .ZN(n97) );
  XOR2_X2 U119 ( .A(n14), .B(n101), .Z(SUM[6]) );
  NAND2_X2 U121 ( .A1(n138), .A2(n100), .ZN(n14) );
  NAND2_X2 U124 ( .A1(A[6]), .A2(B[6]), .ZN(n100) );
  XOR2_X2 U125 ( .A(n15), .B(n106), .Z(SUM[5]) );
  NAND2_X2 U129 ( .A1(n139), .A2(n105), .ZN(n15) );
  NAND2_X2 U132 ( .A1(A[5]), .A2(B[5]), .ZN(n105) );
  XNOR2_X2 U133 ( .A(n111), .B(n16), .ZN(SUM[4]) );
  NAND2_X2 U137 ( .A1(n140), .A2(n110), .ZN(n16) );
  NAND2_X2 U140 ( .A1(A[4]), .A2(B[4]), .ZN(n110) );
  XNOR2_X2 U141 ( .A(n117), .B(n17), .ZN(SUM[3]) );
  NAND2_X2 U146 ( .A1(n141), .A2(n116), .ZN(n17) );
  NAND2_X2 U149 ( .A1(A[3]), .A2(B[3]), .ZN(n116) );
  XOR2_X2 U150 ( .A(n18), .B(n120), .Z(SUM[2]) );
  NAND2_X2 U152 ( .A1(n142), .A2(n119), .ZN(n18) );
  NAND2_X2 U155 ( .A1(A[2]), .A2(B[2]), .ZN(n119) );
  XOR2_X2 U156 ( .A(n124), .B(n19), .Z(SUM[1]) );
  NAND2_X2 U159 ( .A1(n143), .A2(n123), .ZN(n19) );
  NAND2_X2 U162 ( .A1(A[1]), .A2(B[1]), .ZN(n123) );
  XNOR2_X2 U163 ( .A(A[0]), .B(B[0]), .ZN(SUM[0]) );
  AOI21_X2 U168 ( .B1(n111), .B2(n102), .A(n103), .ZN(n101) );
  AOI21_X2 U169 ( .B1(n68), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X2 U170 ( .B1(n91), .B2(n48), .A(n49), .ZN(n47) );
  NOR2_X2 U171 ( .A1(n69), .A2(n50), .ZN(n48) );
  OAI21_X2 U172 ( .B1(n70), .B2(n50), .A(n51), .ZN(n49) );
  OAI21_X2 U173 ( .B1(n90), .B2(n81), .A(n82), .ZN(n80) );
  OAI21_X2 U174 ( .B1(n90), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X2 U175 ( .B1(n46), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X2 U176 ( .B1(n46), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X2 U177 ( .B1(n71), .B2(n84), .A(n72), .ZN(n70) );
  OAI21_X2 U178 ( .B1(n73), .B2(n79), .A(n74), .ZN(n72) );
  AOI21_X2 U179 ( .B1(n211), .B2(n43), .A(n38), .ZN(n36) );
  AOI21_X2 U180 ( .B1(n113), .B2(n121), .A(n114), .ZN(n112) );
  NOR2_X2 U181 ( .A1(n118), .A2(n115), .ZN(n113) );
  OAI21_X2 U182 ( .B1(n115), .B2(n119), .A(n116), .ZN(n114) );
  OAI21_X2 U183 ( .B1(n36), .B2(n30), .A(n31), .ZN(n29) );
  OAI21_X2 U184 ( .B1(n62), .B2(n66), .A(n63), .ZN(n61) );
  OAI21_X2 U185 ( .B1(n104), .B2(n110), .A(n105), .ZN(n103) );
  OAI21_X2 U186 ( .B1(n112), .B2(n92), .A(n93), .ZN(n91) );
  AOI21_X2 U187 ( .B1(n94), .B2(n103), .A(n95), .ZN(n93) );
  NOR2_X2 U188 ( .A1(n99), .A2(n96), .ZN(n94) );
  AOI21_X2 U189 ( .B1(n52), .B2(n61), .A(n53), .ZN(n51) );
  OAI21_X2 U190 ( .B1(n54), .B2(n58), .A(n55), .ZN(n53) );
  AOI21_X2 U191 ( .B1(n29), .B2(n213), .A(n24), .ZN(n22) );
  AOI21_X2 U192 ( .B1(n80), .B2(n76), .A(n77), .ZN(n75) );
  AOI21_X2 U193 ( .B1(n46), .B2(n212), .A(n43), .ZN(n41) );
  OAI21_X2 U194 ( .B1(n122), .B2(n124), .A(n123), .ZN(n121) );
  OAI21_X2 U195 ( .B1(n85), .B2(n89), .A(n86), .ZN(n84) );
  OAI21_X2 U196 ( .B1(n96), .B2(n100), .A(n97), .ZN(n95) );
  OAI21_X2 U197 ( .B1(n101), .B2(n99), .A(n100), .ZN(n98) );
  OAI21_X2 U198 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X2 U199 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  NOR2_X2 U200 ( .A1(n57), .A2(n54), .ZN(n52) );
  NOR2_X2 U201 ( .A1(n78), .A2(n73), .ZN(n71) );
  NOR2_X2 U202 ( .A1(n109), .A2(n104), .ZN(n102) );
  NOR2_X2 U203 ( .A1(n65), .A2(n62), .ZN(n60) );
  NOR2_X2 U204 ( .A1(n35), .A2(n30), .ZN(n28) );
  NOR2_X2 U205 ( .A1(n88), .A2(n85), .ZN(n83) );
  AOI21_X2 U206 ( .B1(n111), .B2(n140), .A(n108), .ZN(n106) );
  OAI21_X2 U207 ( .B1(n120), .B2(n118), .A(n119), .ZN(n117) );
  OAI21_X2 U208 ( .B1(n90), .B2(n88), .A(n89), .ZN(n87) );
  NOR2_X2 U209 ( .A1(A[3]), .A2(B[3]), .ZN(n115) );
  NOR2_X2 U210 ( .A1(A[7]), .A2(B[7]), .ZN(n96) );
  NOR2_X2 U211 ( .A1(A[5]), .A2(B[5]), .ZN(n104) );
  NOR2_X2 U212 ( .A1(A[15]), .A2(B[15]), .ZN(n54) );
  NOR2_X2 U213 ( .A1(A[13]), .A2(B[13]), .ZN(n62) );
  NOR2_X2 U214 ( .A1(A[11]), .A2(B[11]), .ZN(n73) );
  NOR2_X2 U215 ( .A1(A[9]), .A2(B[9]), .ZN(n85) );
  NOR2_X2 U216 ( .A1(A[18]), .A2(B[18]), .ZN(n30) );
  NOR2_X2 U217 ( .A1(A[2]), .A2(B[2]), .ZN(n118) );
  NOR2_X2 U218 ( .A1(A[6]), .A2(B[6]), .ZN(n99) );
  NOR2_X2 U219 ( .A1(A[8]), .A2(B[8]), .ZN(n88) );
  NOR2_X2 U220 ( .A1(A[12]), .A2(B[12]), .ZN(n65) );
  NOR2_X2 U221 ( .A1(A[14]), .A2(B[14]), .ZN(n57) );
  NOR2_X2 U222 ( .A1(A[1]), .A2(B[1]), .ZN(n122) );
  NOR2_X2 U223 ( .A1(A[0]), .A2(B[0]), .ZN(n124) );
  NOR2_X2 U224 ( .A1(A[4]), .A2(B[4]), .ZN(n109) );
  NOR2_X2 U225 ( .A1(A[10]), .A2(B[10]), .ZN(n78) );
  OAI21_X2 U226 ( .B1(n47), .B2(n21), .A(n22), .ZN(CO) );
  OR2_X1 U227 ( .A1(A[17]), .A2(B[17]), .ZN(n211) );
  OR2_X1 U228 ( .A1(A[16]), .A2(B[16]), .ZN(n212) );
  OR2_X1 U229 ( .A1(A[19]), .A2(B[19]), .ZN(n213) );
  INV_X4 U230 ( .A(n91), .ZN(n90) );
  INV_X4 U231 ( .A(n84), .ZN(n82) );
  INV_X4 U232 ( .A(n83), .ZN(n81) );
  INV_X4 U233 ( .A(n79), .ZN(n77) );
  INV_X4 U234 ( .A(n68), .ZN(n67) );
  INV_X4 U235 ( .A(n47), .ZN(n46) );
  INV_X4 U236 ( .A(n45), .ZN(n43) );
  INV_X4 U237 ( .A(n40), .ZN(n38) );
  INV_X4 U238 ( .A(n36), .ZN(n34) );
  INV_X4 U239 ( .A(n35), .ZN(n33) );
  INV_X4 U240 ( .A(n26), .ZN(n24) );
  INV_X4 U241 ( .A(n122), .ZN(n143) );
  INV_X4 U242 ( .A(n118), .ZN(n142) );
  INV_X4 U243 ( .A(n115), .ZN(n141) );
  INV_X4 U244 ( .A(n104), .ZN(n139) );
  INV_X4 U245 ( .A(n99), .ZN(n138) );
  INV_X4 U246 ( .A(n96), .ZN(n137) );
  INV_X4 U247 ( .A(n88), .ZN(n136) );
  INV_X4 U248 ( .A(n85), .ZN(n135) );
  INV_X4 U249 ( .A(n78), .ZN(n76) );
  INV_X4 U250 ( .A(n73), .ZN(n133) );
  INV_X4 U251 ( .A(n65), .ZN(n132) );
  INV_X4 U252 ( .A(n62), .ZN(n131) );
  INV_X4 U253 ( .A(n57), .ZN(n130) );
  INV_X4 U254 ( .A(n54), .ZN(n129) );
  INV_X4 U255 ( .A(n30), .ZN(n126) );
  INV_X4 U256 ( .A(n121), .ZN(n120) );
  INV_X4 U257 ( .A(n112), .ZN(n111) );
  INV_X4 U258 ( .A(n110), .ZN(n108) );
  INV_X4 U259 ( .A(n109), .ZN(n140) );
endmodule


module pipleline_stage_2 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   n105;
  wire   [20:0] stage_result;

  pipleline_stage_2_DW01_add_1 stage_add ( .A(divided[26:7]), .B(divisor), 
        .CI(1'b1), .SUM(stage_result[19:0]), .CO(stage_result[20]) );
  INV_X4 U4 ( .A(1'b1), .ZN(stage_out[0]) );
  INV_X4 U6 ( .A(n105), .ZN(q) );
  BUF_X4 U7 ( .A(divided[0]), .Z(stage_out[1]) );
  BUF_X4 U8 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U9 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U10 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U11 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U12 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U13 ( .A(divided[6]), .Z(stage_out[7]) );
  XNOR2_X2 U14 ( .A(divided[27]), .B(stage_result[20]), .ZN(n105) );
  MUX2_X2 U15 ( .A(divided[7]), .B(stage_result[0]), .S(q), .Z(stage_out[8])
         );
  MUX2_X2 U16 ( .A(divided[8]), .B(stage_result[1]), .S(q), .Z(stage_out[9])
         );
  MUX2_X2 U17 ( .A(divided[9]), .B(stage_result[2]), .S(q), .Z(stage_out[10])
         );
  MUX2_X2 U18 ( .A(divided[10]), .B(stage_result[3]), .S(q), .Z(stage_out[11])
         );
  MUX2_X2 U19 ( .A(divided[11]), .B(stage_result[4]), .S(q), .Z(stage_out[12])
         );
  MUX2_X2 U20 ( .A(divided[12]), .B(stage_result[5]), .S(q), .Z(stage_out[13])
         );
  MUX2_X2 U21 ( .A(divided[13]), .B(stage_result[6]), .S(q), .Z(stage_out[14])
         );
  MUX2_X2 U22 ( .A(divided[14]), .B(stage_result[7]), .S(q), .Z(stage_out[15])
         );
  MUX2_X2 U23 ( .A(divided[15]), .B(stage_result[8]), .S(q), .Z(stage_out[16])
         );
  MUX2_X2 U24 ( .A(divided[16]), .B(stage_result[9]), .S(q), .Z(stage_out[17])
         );
  MUX2_X2 U25 ( .A(divided[17]), .B(stage_result[10]), .S(q), .Z(stage_out[18]) );
  MUX2_X2 U26 ( .A(divided[18]), .B(stage_result[11]), .S(q), .Z(stage_out[19]) );
  MUX2_X2 U27 ( .A(divided[19]), .B(stage_result[12]), .S(q), .Z(stage_out[20]) );
  MUX2_X2 U28 ( .A(divided[20]), .B(stage_result[13]), .S(q), .Z(stage_out[21]) );
  MUX2_X2 U29 ( .A(divided[21]), .B(stage_result[14]), .S(q), .Z(stage_out[22]) );
  MUX2_X2 U30 ( .A(divided[22]), .B(stage_result[15]), .S(q), .Z(stage_out[23]) );
  MUX2_X2 U31 ( .A(divided[23]), .B(stage_result[16]), .S(q), .Z(stage_out[24]) );
  MUX2_X2 U32 ( .A(divided[24]), .B(stage_result[17]), .S(q), .Z(stage_out[25]) );
  MUX2_X2 U33 ( .A(divided[25]), .B(stage_result[18]), .S(q), .Z(stage_out[26]) );
  MUX2_X2 U34 ( .A(divided[26]), .B(stage_result[19]), .S(q), .Z(stage_out[27]) );
endmodule


module pipleline_stage_0 ( divided, divisor, q, stage_out );
  input [27:0] divided;
  input [19:0] divisor;
  output [27:0] stage_out;
  output q;
  wire   \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 ,
         \U4/Z_7 , \U4/Z_8 , \U4/Z_9 , \U4/Z_10 , \U4/Z_11 , \U4/Z_12 ,
         \U4/Z_13 , \U4/Z_14 , \U4/Z_15 , \U4/Z_16 , \U4/Z_17 , \U4/Z_18 ,
         \U4/Z_19 , \U4/DATA2_0 , \U4/DATA2_1 , \U4/DATA2_2 , \U4/DATA2_3 ,
         \U4/DATA2_4 , \U4/DATA2_5 , \U4/DATA2_6 , \U4/DATA2_7 , \U4/DATA2_8 ,
         \U4/DATA2_9 , \U4/DATA2_10 , \U4/DATA2_11 , \U4/DATA2_12 ,
         \U4/DATA2_13 , \U4/DATA2_14 , \U4/DATA2_15 , \U4/DATA2_16 ,
         \U4/DATA2_17 , \U4/DATA2_18 , \U4/DATA2_19 , \stage_add/B[0] ,
         \stage_add/B[1] , \stage_add/B[2] , \stage_add/B[3] ,
         \stage_add/B[4] , \stage_add/B[5] , \stage_add/B[6] ,
         \stage_add/B[7] , \stage_add/B[8] , \stage_add/B[9] ,
         \stage_add/B[10] , \stage_add/B[11] , \stage_add/B[12] ,
         \stage_add/B[13] , \stage_add/B[14] , \stage_add/B[15] ,
         \stage_add/B[16] , \stage_add/B[17] , \stage_add/B[18] ,
         \stage_add/B[19] , n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287;
  assign stage_out[8] = \U4/Z_0 ;
  assign stage_out[9] = \U4/Z_1 ;
  assign stage_out[10] = \U4/Z_2 ;
  assign stage_out[11] = \U4/Z_3 ;
  assign stage_out[12] = \U4/Z_4 ;
  assign stage_out[13] = \U4/Z_5 ;
  assign stage_out[14] = \U4/Z_6 ;
  assign stage_out[15] = \U4/Z_7 ;
  assign stage_out[16] = \U4/Z_8 ;
  assign stage_out[17] = \U4/Z_9 ;
  assign stage_out[18] = \U4/Z_10 ;
  assign stage_out[19] = \U4/Z_11 ;
  assign stage_out[20] = \U4/Z_12 ;
  assign stage_out[21] = \U4/Z_13 ;
  assign stage_out[22] = \U4/Z_14 ;
  assign stage_out[23] = \U4/Z_15 ;
  assign stage_out[24] = \U4/Z_16 ;
  assign stage_out[25] = \U4/Z_17 ;
  assign stage_out[26] = \U4/Z_18 ;
  assign stage_out[27] = \U4/Z_19 ;
  assign \U4/DATA2_0  = divided[7];
  assign \U4/DATA2_1  = divided[8];
  assign \U4/DATA2_2  = divided[9];
  assign \U4/DATA2_3  = divided[10];
  assign \U4/DATA2_4  = divided[11];
  assign \U4/DATA2_5  = divided[12];
  assign \U4/DATA2_6  = divided[13];
  assign \U4/DATA2_7  = divided[14];
  assign \U4/DATA2_8  = divided[15];
  assign \U4/DATA2_9  = divided[16];
  assign \U4/DATA2_10  = divided[17];
  assign \U4/DATA2_11  = divided[18];
  assign \U4/DATA2_12  = divided[19];
  assign \U4/DATA2_13  = divided[20];
  assign \U4/DATA2_14  = divided[21];
  assign \U4/DATA2_15  = divided[22];
  assign \U4/DATA2_16  = divided[23];
  assign \U4/DATA2_17  = divided[24];
  assign \U4/DATA2_18  = divided[25];
  assign \U4/DATA2_19  = divided[26];
  assign \stage_add/B[0]  = divisor[0];
  assign \stage_add/B[1]  = divisor[1];
  assign \stage_add/B[2]  = divisor[2];
  assign \stage_add/B[3]  = divisor[3];
  assign \stage_add/B[4]  = divisor[4];
  assign \stage_add/B[5]  = divisor[5];
  assign \stage_add/B[6]  = divisor[6];
  assign \stage_add/B[7]  = divisor[7];
  assign \stage_add/B[8]  = divisor[8];
  assign \stage_add/B[9]  = divisor[9];
  assign \stage_add/B[10]  = divisor[10];
  assign \stage_add/B[11]  = divisor[11];
  assign \stage_add/B[12]  = divisor[12];
  assign \stage_add/B[13]  = divisor[13];
  assign \stage_add/B[14]  = divisor[14];
  assign \stage_add/B[15]  = divisor[15];
  assign \stage_add/B[16]  = divisor[16];
  assign \stage_add/B[17]  = divisor[17];
  assign \stage_add/B[18]  = divisor[18];
  assign \stage_add/B[19]  = divisor[19];

  INV_X4 U3 ( .A(1'b1), .ZN(stage_out[0]) );
  AND3_X2 U5 ( .A1(n121), .A2(n122), .A3(n259), .ZN(n125) );
  NAND2_X2 U6 ( .A1(n164), .A2(n165), .ZN(n277) );
  OR2_X4 U7 ( .A1(n183), .A2(n182), .ZN(n98) );
  NOR2_X4 U8 ( .A1(n153), .A2(n103), .ZN(n158) );
  NAND2_X2 U9 ( .A1(n118), .A2(n119), .ZN(n120) );
  OAI21_X2 U10 ( .B1(\stage_add/B[10] ), .B2(\U4/DATA2_10 ), .A(n234), .ZN(
        n240) );
  NAND3_X2 U11 ( .A1(n171), .A2(n102), .A3(n179), .ZN(n177) );
  NAND2_X2 U12 ( .A1(n184), .A2(n143), .ZN(n186) );
  OAI211_X4 U13 ( .C1(n158), .C2(n157), .A(n156), .B(n247), .ZN(n253) );
  AND2_X4 U14 ( .A1(n206), .A2(n210), .ZN(n99) );
  AND2_X4 U15 ( .A1(n230), .A2(n236), .ZN(n100) );
  AND2_X4 U16 ( .A1(n99), .A2(n104), .ZN(n101) );
  NAND2_X2 U17 ( .A1(n109), .A2(n110), .ZN(n102) );
  OR2_X4 U18 ( .A1(n227), .A2(n240), .ZN(n103) );
  AND2_X4 U19 ( .A1(n192), .A2(n198), .ZN(n104) );
  AND2_X4 U20 ( .A1(n223), .A2(n217), .ZN(n105) );
  AND2_X4 U21 ( .A1(n178), .A2(n172), .ZN(n106) );
  NAND2_X2 U22 ( .A1(n106), .A2(n117), .ZN(n176) );
  AND2_X4 U23 ( .A1(n99), .A2(n202), .ZN(n107) );
  AND2_X1 U24 ( .A1(n142), .A2(n141), .ZN(n108) );
  NOR3_X1 U25 ( .A1(n107), .A2(n108), .A3(n131), .ZN(n148) );
  NAND2_X1 U26 ( .A1(n277), .A2(n112), .ZN(n109) );
  OR2_X1 U27 ( .A1(n111), .A2(n167), .ZN(n110) );
  INV_X4 U28 ( .A(n168), .ZN(n111) );
  AND2_X1 U29 ( .A1(n116), .A2(n168), .ZN(n112) );
  NOR2_X4 U30 ( .A1(n183), .A2(n182), .ZN(n113) );
  INV_X4 U31 ( .A(n98), .ZN(n114) );
  INV_X4 U32 ( .A(n113), .ZN(q) );
  NAND2_X1 U33 ( .A1(n275), .A2(q), .ZN(n276) );
  NAND2_X1 U34 ( .A1(n263), .A2(n98), .ZN(n264) );
  NAND2_X1 U35 ( .A1(n251), .A2(q), .ZN(n252) );
  NAND2_X1 U36 ( .A1(n238), .A2(n98), .ZN(n239) );
  NAND2_X1 U37 ( .A1(n225), .A2(q), .ZN(n226) );
  NAND2_X1 U38 ( .A1(n200), .A2(n98), .ZN(n201) );
  INV_X1 U39 ( .A(n117), .ZN(n284) );
  NAND2_X2 U40 ( .A1(n101), .A2(n203), .ZN(n147) );
  OR2_X1 U41 ( .A1(\stage_add/B[17] ), .A2(\U4/DATA2_17 ), .ZN(n116) );
  NAND2_X2 U42 ( .A1(n116), .A2(n277), .ZN(n166) );
  NAND2_X1 U43 ( .A1(n217), .A2(n216), .ZN(n220) );
  INV_X2 U44 ( .A(\stage_add/B[3] ), .ZN(n139) );
  NAND2_X1 U45 ( .A1(n104), .A2(n203), .ZN(n204) );
  NAND2_X1 U46 ( .A1(n192), .A2(n203), .ZN(n195) );
  OAI22_X1 U47 ( .A1(n185), .A2(n184), .B1(n114), .B2(n186), .ZN(\U4/Z_0 ) );
  INV_X2 U48 ( .A(n186), .ZN(n124) );
  NAND2_X1 U49 ( .A1(\stage_add/B[2] ), .A2(\U4/DATA2_2 ), .ZN(n192) );
  BUF_X4 U50 ( .A(divided[6]), .Z(stage_out[7]) );
  BUF_X4 U51 ( .A(divided[5]), .Z(stage_out[6]) );
  BUF_X4 U52 ( .A(divided[4]), .Z(stage_out[5]) );
  BUF_X4 U53 ( .A(divided[3]), .Z(stage_out[4]) );
  BUF_X4 U54 ( .A(divided[2]), .Z(stage_out[3]) );
  BUF_X4 U55 ( .A(divided[1]), .Z(stage_out[2]) );
  BUF_X4 U56 ( .A(divided[0]), .Z(stage_out[1]) );
  NAND2_X2 U57 ( .A1(n168), .A2(n280), .ZN(n117) );
  NAND2_X2 U58 ( .A1(n105), .A2(n216), .ZN(n228) );
  NAND2_X1 U59 ( .A1(\stage_add/B[6] ), .A2(\U4/DATA2_6 ), .ZN(n217) );
  NAND2_X1 U60 ( .A1(\stage_add/B[7] ), .A2(\U4/DATA2_7 ), .ZN(n223) );
  NAND2_X1 U61 ( .A1(n229), .A2(n228), .ZN(n241) );
  NAND2_X2 U62 ( .A1(n120), .A2(n196), .ZN(n202) );
  INV_X1 U63 ( .A(\stage_add/B[4] ), .ZN(n118) );
  INV_X1 U64 ( .A(\U4/DATA2_4 ), .ZN(n119) );
  OR2_X4 U65 ( .A1(n123), .A2(n124), .ZN(n144) );
  OAI21_X2 U66 ( .B1(\stage_add/B[8] ), .B2(\U4/DATA2_8 ), .A(n221), .ZN(n227)
         );
  NAND2_X2 U67 ( .A1(n126), .A2(n127), .ZN(n121) );
  NAND2_X2 U68 ( .A1(n253), .A2(n128), .ZN(n122) );
  INV_X4 U69 ( .A(\stage_add/B[14] ), .ZN(n126) );
  INV_X4 U70 ( .A(\U4/DATA2_14 ), .ZN(n127) );
  INV_X1 U71 ( .A(n125), .ZN(n265) );
  NOR2_X1 U72 ( .A1(\U4/DATA2_5 ), .A2(\stage_add/B[5] ), .ZN(n131) );
  NOR2_X2 U73 ( .A1(\stage_add/B[1] ), .A2(\U4/DATA2_1 ), .ZN(n123) );
  AND2_X4 U74 ( .A1(n254), .A2(n261), .ZN(n128) );
  XOR2_X1 U75 ( .A(\U4/DATA2_3 ), .B(n194), .Z(\U4/Z_3 ) );
  XOR2_X1 U76 ( .A(\U4/DATA2_6 ), .B(n215), .Z(\U4/Z_6 ) );
  XOR2_X1 U77 ( .A(\U4/DATA2_7 ), .B(n219), .Z(\U4/Z_7 ) );
  XOR2_X1 U78 ( .A(\U4/DATA2_9 ), .B(n232), .Z(\U4/Z_9 ) );
  XOR2_X1 U79 ( .A(\U4/DATA2_1 ), .B(n188), .Z(\U4/Z_1 ) );
  XOR2_X1 U80 ( .A(\U4/DATA2_5 ), .B(n209), .Z(\U4/Z_5 ) );
  XOR2_X1 U81 ( .A(\U4/DATA2_2 ), .B(n191), .Z(\U4/Z_2 ) );
  XOR2_X1 U82 ( .A(\U4/DATA2_11 ), .B(n245), .Z(\U4/Z_11 ) );
  XNOR2_X1 U83 ( .A(\U4/DATA2_4 ), .B(n201), .ZN(\U4/Z_4 ) );
  XNOR2_X1 U84 ( .A(\U4/DATA2_8 ), .B(n226), .ZN(\U4/Z_8 ) );
  XNOR2_X1 U85 ( .A(\U4/DATA2_10 ), .B(n239), .ZN(\U4/Z_10 ) );
  INV_X1 U86 ( .A(n202), .ZN(n205) );
  OR2_X2 U87 ( .A1(\U4/DATA2_11 ), .A2(\stage_add/B[11] ), .ZN(n247) );
  XNOR2_X1 U88 ( .A(\stage_add/B[1] ), .B(n186), .ZN(n187) );
  XNOR2_X1 U89 ( .A(\stage_add/B[2] ), .B(n189), .ZN(n190) );
  XNOR2_X1 U90 ( .A(\stage_add/B[3] ), .B(n195), .ZN(n193) );
  XNOR2_X1 U91 ( .A(\stage_add/B[7] ), .B(n220), .ZN(n218) );
  XNOR2_X1 U92 ( .A(\stage_add/B[9] ), .B(n233), .ZN(n231) );
  XNOR2_X1 U93 ( .A(\stage_add/B[11] ), .B(n246), .ZN(n244) );
  XNOR2_X1 U94 ( .A(\stage_add/B[17] ), .B(n277), .ZN(n278) );
  XNOR2_X1 U95 ( .A(\stage_add/B[18] ), .B(n280), .ZN(n281) );
  XOR2_X1 U96 ( .A(n199), .B(\stage_add/B[4] ), .Z(n200) );
  NAND2_X1 U97 ( .A1(n198), .A2(n197), .ZN(n199) );
  XOR2_X1 U98 ( .A(n224), .B(\stage_add/B[8] ), .Z(n225) );
  NAND2_X1 U99 ( .A1(n223), .A2(n222), .ZN(n224) );
  XOR2_X1 U100 ( .A(n237), .B(\stage_add/B[10] ), .Z(n238) );
  NAND2_X1 U101 ( .A1(n236), .A2(n235), .ZN(n237) );
  NAND2_X1 U102 ( .A1(n249), .A2(n248), .ZN(n250) );
  OAI211_X2 U103 ( .C1(n100), .C2(n240), .A(n249), .B(n242), .ZN(n157) );
  OR2_X1 U104 ( .A1(n240), .A2(n129), .ZN(n243) );
  AND2_X4 U105 ( .A1(n100), .A2(n241), .ZN(n129) );
  AND2_X1 U106 ( .A1(n207), .A2(n206), .ZN(n130) );
  OR2_X1 U107 ( .A1(\U4/DATA2_18 ), .A2(\stage_add/B[18] ), .ZN(n168) );
  OR2_X1 U108 ( .A1(\U4/DATA2_2 ), .A2(\stage_add/B[2] ), .ZN(n146) );
  XOR2_X2 U109 ( .A(n250), .B(\stage_add/B[12] ), .Z(n251) );
  XOR2_X2 U110 ( .A(n262), .B(\stage_add/B[14] ), .Z(n263) );
  XOR2_X2 U111 ( .A(n274), .B(\stage_add/B[16] ), .Z(n275) );
  INV_X4 U112 ( .A(divided[27]), .ZN(n171) );
  NAND2_X2 U113 ( .A1(\U4/DATA2_17 ), .A2(\stage_add/B[17] ), .ZN(n167) );
  NAND2_X2 U114 ( .A1(\stage_add/B[16] ), .A2(\U4/DATA2_16 ), .ZN(n165) );
  NAND2_X2 U115 ( .A1(\stage_add/B[4] ), .A2(\U4/DATA2_4 ), .ZN(n206) );
  NAND2_X2 U116 ( .A1(\stage_add/B[5] ), .A2(\U4/DATA2_5 ), .ZN(n210) );
  INV_X4 U117 ( .A(\U4/DATA2_3 ), .ZN(n140) );
  NAND2_X2 U118 ( .A1(n140), .A2(n139), .ZN(n196) );
  INV_X4 U119 ( .A(\U4/DATA2_6 ), .ZN(n142) );
  INV_X4 U120 ( .A(\stage_add/B[6] ), .ZN(n141) );
  NAND2_X2 U121 ( .A1(\stage_add/B[3] ), .A2(\U4/DATA2_3 ), .ZN(n198) );
  NAND2_X2 U122 ( .A1(\U4/DATA2_1 ), .A2(\stage_add/B[1] ), .ZN(n145) );
  INV_X4 U123 ( .A(\U4/DATA2_0 ), .ZN(n184) );
  INV_X4 U124 ( .A(\stage_add/B[0] ), .ZN(n143) );
  NAND2_X2 U125 ( .A1(n145), .A2(n144), .ZN(n189) );
  NAND2_X2 U126 ( .A1(n189), .A2(n146), .ZN(n203) );
  NAND2_X2 U127 ( .A1(n148), .A2(n147), .ZN(n216) );
  INV_X4 U128 ( .A(n228), .ZN(n153) );
  INV_X4 U129 ( .A(\U4/DATA2_9 ), .ZN(n150) );
  INV_X4 U130 ( .A(\stage_add/B[9] ), .ZN(n149) );
  NAND2_X2 U131 ( .A1(n150), .A2(n149), .ZN(n234) );
  INV_X4 U132 ( .A(\U4/DATA2_7 ), .ZN(n152) );
  INV_X4 U133 ( .A(\stage_add/B[7] ), .ZN(n151) );
  NAND2_X2 U134 ( .A1(n152), .A2(n151), .ZN(n221) );
  NAND2_X2 U135 ( .A1(\stage_add/B[8] ), .A2(\U4/DATA2_8 ), .ZN(n230) );
  NAND2_X2 U136 ( .A1(\stage_add/B[9] ), .A2(\U4/DATA2_9 ), .ZN(n236) );
  NAND2_X2 U137 ( .A1(\stage_add/B[11] ), .A2(\U4/DATA2_11 ), .ZN(n249) );
  NAND2_X2 U138 ( .A1(\stage_add/B[10] ), .A2(\U4/DATA2_10 ), .ZN(n242) );
  INV_X4 U139 ( .A(\U4/DATA2_12 ), .ZN(n155) );
  INV_X4 U140 ( .A(\stage_add/B[12] ), .ZN(n154) );
  NAND2_X2 U141 ( .A1(n155), .A2(n154), .ZN(n156) );
  NAND2_X2 U142 ( .A1(\stage_add/B[12] ), .A2(\U4/DATA2_12 ), .ZN(n254) );
  NAND2_X2 U143 ( .A1(\stage_add/B[13] ), .A2(\U4/DATA2_13 ), .ZN(n261) );
  INV_X4 U144 ( .A(\U4/DATA2_13 ), .ZN(n160) );
  INV_X4 U145 ( .A(\stage_add/B[13] ), .ZN(n159) );
  NAND2_X2 U146 ( .A1(n160), .A2(n159), .ZN(n259) );
  NAND2_X2 U147 ( .A1(\stage_add/B[14] ), .A2(\U4/DATA2_14 ), .ZN(n266) );
  NAND2_X2 U148 ( .A1(\stage_add/B[15] ), .A2(\U4/DATA2_15 ), .ZN(n273) );
  NAND2_X2 U149 ( .A1(n266), .A2(n273), .ZN(n163) );
  INV_X4 U150 ( .A(\U4/DATA2_15 ), .ZN(n162) );
  INV_X4 U151 ( .A(\stage_add/B[15] ), .ZN(n161) );
  NAND2_X2 U152 ( .A1(n162), .A2(n161), .ZN(n271) );
  OAI221_X2 U153 ( .B1(\stage_add/B[16] ), .B2(\U4/DATA2_16 ), .C1(n125), .C2(
        n163), .A(n271), .ZN(n164) );
  NAND2_X2 U154 ( .A1(n167), .A2(n166), .ZN(n280) );
  INV_X4 U155 ( .A(\U4/DATA2_19 ), .ZN(n170) );
  INV_X4 U156 ( .A(\stage_add/B[19] ), .ZN(n169) );
  NAND2_X2 U157 ( .A1(n170), .A2(n169), .ZN(n179) );
  NAND2_X2 U158 ( .A1(\stage_add/B[18] ), .A2(\U4/DATA2_18 ), .ZN(n178) );
  NAND2_X2 U159 ( .A1(\stage_add/B[19] ), .A2(\U4/DATA2_19 ), .ZN(n173) );
  NAND2_X2 U160 ( .A1(divided[27]), .A2(n173), .ZN(n180) );
  INV_X4 U161 ( .A(n180), .ZN(n172) );
  INV_X4 U162 ( .A(n173), .ZN(n174) );
  NAND2_X2 U163 ( .A1(n174), .A2(n171), .ZN(n175) );
  NAND3_X2 U164 ( .A1(n177), .A2(n176), .A3(n175), .ZN(n183) );
  INV_X4 U165 ( .A(n178), .ZN(n283) );
  NAND2_X2 U166 ( .A1(n283), .A2(n179), .ZN(n181) );
  OAI22_X2 U167 ( .A1(divided[27]), .A2(n181), .B1(n180), .B2(n179), .ZN(n182)
         );
  NOR2_X2 U168 ( .A1(\stage_add/B[0] ), .A2(n114), .ZN(n185) );
  NOR2_X2 U169 ( .A1(n114), .A2(n187), .ZN(n188) );
  NOR2_X2 U170 ( .A1(n114), .A2(n190), .ZN(n191) );
  NOR2_X2 U171 ( .A1(n114), .A2(n193), .ZN(n194) );
  NAND2_X2 U172 ( .A1(n196), .A2(n195), .ZN(n197) );
  NAND2_X2 U173 ( .A1(n205), .A2(n204), .ZN(n207) );
  XOR2_X2 U174 ( .A(\stage_add/B[5] ), .B(n130), .Z(n208) );
  NOR2_X2 U175 ( .A1(n114), .A2(n208), .ZN(n209) );
  INV_X4 U176 ( .A(n210), .ZN(n212) );
  NOR2_X2 U177 ( .A1(n131), .A2(n130), .ZN(n211) );
  NOR2_X2 U178 ( .A1(n212), .A2(n211), .ZN(n213) );
  XOR2_X2 U179 ( .A(\stage_add/B[6] ), .B(n213), .Z(n214) );
  NOR2_X2 U180 ( .A1(n114), .A2(n214), .ZN(n215) );
  NOR2_X2 U181 ( .A1(n114), .A2(n218), .ZN(n219) );
  NAND2_X2 U182 ( .A1(n221), .A2(n220), .ZN(n222) );
  INV_X4 U183 ( .A(n227), .ZN(n229) );
  NAND2_X2 U184 ( .A1(n241), .A2(n230), .ZN(n233) );
  NOR2_X2 U185 ( .A1(n114), .A2(n231), .ZN(n232) );
  NAND2_X2 U186 ( .A1(n234), .A2(n233), .ZN(n235) );
  NAND2_X2 U187 ( .A1(n243), .A2(n242), .ZN(n246) );
  NOR2_X2 U188 ( .A1(n114), .A2(n244), .ZN(n245) );
  NAND2_X2 U189 ( .A1(n247), .A2(n246), .ZN(n248) );
  XNOR2_X2 U190 ( .A(\U4/DATA2_12 ), .B(n252), .ZN(\U4/Z_12 ) );
  NAND2_X2 U191 ( .A1(n254), .A2(n253), .ZN(n258) );
  INV_X4 U192 ( .A(n258), .ZN(n255) );
  XOR2_X2 U193 ( .A(\stage_add/B[13] ), .B(n255), .Z(n256) );
  NOR2_X2 U194 ( .A1(n114), .A2(n256), .ZN(n257) );
  XOR2_X2 U195 ( .A(\U4/DATA2_13 ), .B(n257), .Z(\U4/Z_13 ) );
  NAND2_X2 U196 ( .A1(n259), .A2(n258), .ZN(n260) );
  NAND2_X2 U197 ( .A1(n261), .A2(n260), .ZN(n262) );
  XNOR2_X2 U198 ( .A(\U4/DATA2_14 ), .B(n264), .ZN(\U4/Z_14 ) );
  NAND2_X2 U199 ( .A1(n266), .A2(n265), .ZN(n270) );
  INV_X4 U200 ( .A(n270), .ZN(n267) );
  XOR2_X2 U201 ( .A(\stage_add/B[15] ), .B(n267), .Z(n268) );
  NOR2_X2 U202 ( .A1(n114), .A2(n268), .ZN(n269) );
  XOR2_X2 U203 ( .A(\U4/DATA2_15 ), .B(n269), .Z(\U4/Z_15 ) );
  NAND2_X2 U204 ( .A1(n271), .A2(n270), .ZN(n272) );
  NAND2_X2 U205 ( .A1(n273), .A2(n272), .ZN(n274) );
  XNOR2_X2 U206 ( .A(\U4/DATA2_16 ), .B(n276), .ZN(\U4/Z_16 ) );
  NOR2_X2 U207 ( .A1(n114), .A2(n278), .ZN(n279) );
  XOR2_X2 U208 ( .A(\U4/DATA2_17 ), .B(n279), .Z(\U4/Z_17 ) );
  NOR2_X2 U209 ( .A1(n114), .A2(n281), .ZN(n282) );
  XOR2_X2 U210 ( .A(\U4/DATA2_18 ), .B(n282), .Z(\U4/Z_18 ) );
  NOR2_X2 U211 ( .A1(n284), .A2(n283), .ZN(n285) );
  XOR2_X2 U212 ( .A(\stage_add/B[19] ), .B(n285), .Z(n286) );
  NOR2_X2 U213 ( .A1(n114), .A2(n286), .ZN(n287) );
  XOR2_X2 U214 ( .A(\U4/DATA2_19 ), .B(n287), .Z(\U4/Z_19 ) );
endmodule


module pipeline_divider ( clock, reset_n, start, divided, divisor, q, StartOut
 );
  input [27:0] divided;
  input [19:0] divisor;
  output [7:0] q;
  input clock, reset_n, start;
  output StartOut;
  wire   n132, n131, n130, n129, n128, n127, n126, n125, n124, n123, n122,
         n121, n120, n119, n118, n117, n116, n115, n114, n113, n160, n159,
         n158, n157, n156, n155, n154, n153, n152, n151, n150, n149, n148,
         n147, n146, n145, n144, n143, n142, n141, n140, n139, n138, n137,
         n136, n135, n134, n245, n299, n298, n297, n296, n295, n294, n293,
         n292, n291, n290, n289, n288, n287, n286, n285, n284, n283, n282,
         n281, n280, n279, n278, n277, n276, n275, n274, n273, n383, n436,
         n435, n434, n433, n432, n431, n430, n429, n428, n427, n426, n425,
         n424, n423, n422, n421, n420, n419, n418, n417, n416, n415, n414,
         n413, n412, n411, n410, n519, n571, n570, n569, n568, n567, n566,
         n565, n564, n563, n562, n561, n560, n559, n558, n557, n556, n555,
         n554, n553, n552, n551, n550, n549, n548, n547, n546, n545, n653,
         n704, n703, n702, n701, n700, n699, n698, n697, n696, n695, n694,
         n693, n692, n691, n690, n689, n688, n687, n686, n685, n684, n683,
         n682, n681, n680, n679, n678, n835, n834, n833, n832, n831, n830,
         n829, n828, n827, n826, n825, n824, n823, n822, n821, n820, n819,
         n818, n817, n816, n815, n814, n813, n812, n811, n810, n809, n915,
         n964, n963, n962, n961, n960, n959, n958, n957, n956, n955, n954,
         n953, n952, n951, n950, n949, n948, n947, n946, n945, n944, n943,
         n942, n941, n940, n939, n938, \U25/Z_1 , \U25/Z_2 , \U25/Z_3 ,
         \U25/Z_4 , \U25/Z_5 , \U25/Z_6 , \U25/Z_7 , \U25/Z_8 , \U25/Z_9 ,
         \U25/Z_10 , \U25/Z_11 , \U25/Z_12 , \U25/Z_13 , \U25/Z_14 ,
         \U25/Z_15 , \U25/Z_16 , \U25/Z_17 , \U25/Z_18 , \U25/Z_19 ,
         \U25/Z_20 , \U25/Z_21 , \U25/Z_22 , \U25/Z_23 , \U25/Z_24 ,
         \U25/Z_25 , \U25/Z_26 , \U25/Z_27 , \U25/DATA1_1 , \U25/DATA1_2 ,
         \U25/DATA1_3 , \U25/DATA1_4 , \U25/DATA1_5 , \U25/DATA1_6 ,
         \U25/DATA1_7 , \U25/DATA1_8 , \U25/DATA1_9 , \U25/DATA1_10 ,
         \U25/DATA1_11 , \U25/DATA1_12 , \U25/DATA1_13 , \U25/DATA1_14 ,
         \U25/DATA1_15 , \U25/DATA1_16 , \U25/DATA1_17 , \U25/DATA1_18 ,
         \U25/DATA1_19 , \U25/DATA1_20 , \U25/DATA1_21 , \U25/DATA1_22 ,
         \U25/DATA1_23 , \U25/DATA1_24 , \U25/DATA1_25 , \U25/DATA1_26 ,
         \U25/DATA1_27 , \U23/Z_0 , \U23/DATA1_0 , \U22/Z_1 , \U22/Z_2 ,
         \U22/Z_3 , \U22/Z_4 , \U22/Z_5 , \U22/Z_6 , \U22/Z_7 , \U22/Z_8 ,
         \U22/Z_9 , \U22/Z_10 , \U22/Z_11 , \U22/Z_12 , \U22/Z_13 , \U22/Z_14 ,
         \U22/Z_15 , \U22/Z_16 , \U22/Z_17 , \U22/Z_18 , \U22/Z_19 ,
         \U22/Z_20 , \U22/Z_21 , \U22/Z_22 , \U22/Z_23 , \U22/Z_24 ,
         \U22/Z_25 , \U22/Z_26 , \U22/Z_27 , \U22/DATA1_1 , \U22/DATA1_2 ,
         \U22/DATA1_3 , \U22/DATA1_4 , \U22/DATA1_5 , \U22/DATA1_6 ,
         \U22/DATA1_7 , \U22/DATA1_8 , \U22/DATA1_9 , \U22/DATA1_10 ,
         \U22/DATA1_11 , \U22/DATA1_12 , \U22/DATA1_13 , \U22/DATA1_14 ,
         \U22/DATA1_15 , \U22/DATA1_16 , \U22/DATA1_17 , \U22/DATA1_18 ,
         \U22/DATA1_19 , \U22/DATA1_20 , \U22/DATA1_21 , \U22/DATA1_22 ,
         \U22/DATA1_23 , \U22/DATA1_24 , \U22/DATA1_25 , \U22/DATA1_26 ,
         \U22/DATA1_27 , \U21/Z_0 , \U21/Z_1 , \U21/Z_2 , \U21/Z_3 , \U21/Z_4 ,
         \U21/Z_5 , \U21/Z_6 , \U21/Z_7 , \U21/Z_8 , \U21/Z_9 , \U21/Z_10 ,
         \U21/Z_11 , \U21/Z_12 , \U21/Z_13 , \U21/Z_14 , \U21/Z_15 ,
         \U21/Z_16 , \U21/Z_17 , \U21/Z_18 , \U21/Z_19 , \U21/DATA1_0 ,
         \U21/DATA1_1 , \U21/DATA1_2 , \U21/DATA1_3 , \U21/DATA1_4 ,
         \U21/DATA1_5 , \U21/DATA1_6 , \U21/DATA1_7 , \U21/DATA1_8 ,
         \U21/DATA1_9 , \U21/DATA1_10 , \U21/DATA1_11 , \U21/DATA1_12 ,
         \U21/DATA1_13 , \U21/DATA1_14 , \U21/DATA1_15 , \U21/DATA1_16 ,
         \U21/DATA1_17 , \U21/DATA1_18 , \U21/DATA1_19 , \U20/Z_0 , \U20/Z_1 ,
         \U20/DATA1_0 , \U20/DATA1_1 , \U19/Z_1 , \U19/Z_2 , \U19/Z_3 ,
         \U19/Z_4 , \U19/Z_5 , \U19/Z_6 , \U19/Z_7 , \U19/Z_8 , \U19/Z_9 ,
         \U19/Z_10 , \U19/Z_11 , \U19/Z_12 , \U19/Z_13 , \U19/Z_14 ,
         \U19/Z_15 , \U19/Z_16 , \U19/Z_17 , \U19/Z_18 , \U19/Z_19 ,
         \U19/Z_20 , \U19/Z_21 , \U19/Z_22 , \U19/Z_23 , \U19/Z_24 ,
         \U19/Z_25 , \U19/Z_26 , \U19/Z_27 , \U19/DATA1_1 , \U19/DATA1_2 ,
         \U19/DATA1_3 , \U19/DATA1_4 , \U19/DATA1_5 , \U19/DATA1_6 ,
         \U19/DATA1_7 , \U19/DATA1_8 , \U19/DATA1_9 , \U19/DATA1_10 ,
         \U19/DATA1_11 , \U19/DATA1_12 , \U19/DATA1_13 , \U19/DATA1_14 ,
         \U19/DATA1_15 , \U19/DATA1_16 , \U19/DATA1_17 , \U19/DATA1_18 ,
         \U19/DATA1_19 , \U19/DATA1_20 , \U19/DATA1_21 , \U19/DATA1_22 ,
         \U19/DATA1_23 , \U19/DATA1_24 , \U19/DATA1_25 , \U19/DATA1_26 ,
         \U19/DATA1_27 , \U18/Z_0 , \U18/Z_1 , \U18/Z_2 , \U18/Z_3 , \U18/Z_4 ,
         \U18/Z_5 , \U18/Z_6 , \U18/Z_7 , \U18/Z_8 , \U18/Z_9 , \U18/Z_10 ,
         \U18/Z_11 , \U18/Z_12 , \U18/Z_13 , \U18/Z_14 , \U18/Z_15 ,
         \U18/Z_16 , \U18/Z_17 , \U18/Z_18 , \U18/Z_19 , \U18/DATA1_0 ,
         \U18/DATA1_1 , \U18/DATA1_2 , \U18/DATA1_3 , \U18/DATA1_4 ,
         \U18/DATA1_5 , \U18/DATA1_6 , \U18/DATA1_7 , \U18/DATA1_8 ,
         \U18/DATA1_9 , \U18/DATA1_10 , \U18/DATA1_11 , \U18/DATA1_12 ,
         \U18/DATA1_13 , \U18/DATA1_14 , \U18/DATA1_15 , \U18/DATA1_16 ,
         \U18/DATA1_17 , \U18/DATA1_18 , \U18/DATA1_19 , \U17/Z_0 , \U17/Z_1 ,
         \U17/Z_2 , \U17/DATA1_0 , \U17/DATA1_1 , \U17/DATA1_2 , \U16/Z_1 ,
         \U16/Z_2 , \U16/Z_3 , \U16/Z_4 , \U16/Z_5 , \U16/Z_6 , \U16/Z_7 ,
         \U16/Z_8 , \U16/Z_9 , \U16/Z_10 , \U16/Z_11 , \U16/Z_12 , \U16/Z_13 ,
         \U16/Z_14 , \U16/Z_15 , \U16/Z_16 , \U16/Z_17 , \U16/Z_18 ,
         \U16/Z_19 , \U16/Z_20 , \U16/Z_21 , \U16/Z_22 , \U16/Z_23 ,
         \U16/Z_24 , \U16/Z_25 , \U16/Z_26 , \U16/Z_27 , \U16/DATA1_1 ,
         \U16/DATA1_2 , \U16/DATA1_3 , \U16/DATA1_4 , \U16/DATA1_5 ,
         \U16/DATA1_6 , \U16/DATA1_7 , \U16/DATA1_8 , \U16/DATA1_9 ,
         \U16/DATA1_10 , \U16/DATA1_11 , \U16/DATA1_12 , \U16/DATA1_13 ,
         \U16/DATA1_14 , \U16/DATA1_15 , \U16/DATA1_16 , \U16/DATA1_17 ,
         \U16/DATA1_18 , \U16/DATA1_19 , \U16/DATA1_20 , \U16/DATA1_21 ,
         \U16/DATA1_22 , \U16/DATA1_23 , \U16/DATA1_24 , \U16/DATA1_25 ,
         \U16/DATA1_26 , \U16/DATA1_27 , \U15/Z_0 , \U15/Z_1 , \U15/Z_2 ,
         \U15/Z_3 , \U15/Z_4 , \U15/Z_5 , \U15/Z_6 , \U15/Z_7 , \U15/Z_8 ,
         \U15/Z_9 , \U15/Z_10 , \U15/Z_11 , \U15/Z_12 , \U15/Z_13 , \U15/Z_14 ,
         \U15/Z_15 , \U15/Z_16 , \U15/Z_17 , \U15/Z_18 , \U15/Z_19 ,
         \U15/DATA1_0 , \U15/DATA1_1 , \U15/DATA1_2 , \U15/DATA1_3 ,
         \U15/DATA1_4 , \U15/DATA1_5 , \U15/DATA1_6 , \U15/DATA1_7 ,
         \U15/DATA1_8 , \U15/DATA1_9 , \U15/DATA1_10 , \U15/DATA1_11 ,
         \U15/DATA1_12 , \U15/DATA1_13 , \U15/DATA1_14 , \U15/DATA1_15 ,
         \U15/DATA1_16 , \U15/DATA1_17 , \U15/DATA1_18 , \U15/DATA1_19 ,
         \U14/Z_0 , \U14/Z_1 , \U14/Z_2 , \U14/Z_3 , \U14/DATA1_0 ,
         \U14/DATA1_1 , \U14/DATA1_2 , \U14/DATA1_3 , \U13/Z_1 , \U13/Z_2 ,
         \U13/Z_3 , \U13/Z_4 , \U13/Z_5 , \U13/Z_6 , \U13/Z_7 , \U13/Z_8 ,
         \U13/Z_9 , \U13/Z_10 , \U13/Z_11 , \U13/Z_12 , \U13/Z_13 , \U13/Z_14 ,
         \U13/Z_15 , \U13/Z_16 , \U13/Z_17 , \U13/Z_18 , \U13/Z_19 ,
         \U13/Z_20 , \U13/Z_21 , \U13/Z_22 , \U13/Z_23 , \U13/Z_24 ,
         \U13/Z_25 , \U13/Z_26 , \U13/Z_27 , \U13/DATA1_1 , \U13/DATA1_2 ,
         \U13/DATA1_3 , \U13/DATA1_4 , \U13/DATA1_5 , \U13/DATA1_6 ,
         \U13/DATA1_7 , \U13/DATA1_8 , \U13/DATA1_9 , \U13/DATA1_10 ,
         \U13/DATA1_11 , \U13/DATA1_12 , \U13/DATA1_13 , \U13/DATA1_14 ,
         \U13/DATA1_15 , \U13/DATA1_16 , \U13/DATA1_17 , \U13/DATA1_18 ,
         \U13/DATA1_19 , \U13/DATA1_20 , \U13/DATA1_21 , \U13/DATA1_22 ,
         \U13/DATA1_23 , \U13/DATA1_24 , \U13/DATA1_25 , \U13/DATA1_26 ,
         \U13/DATA1_27 , \U12/Z_0 , \U12/Z_1 , \U12/Z_2 , \U12/Z_3 , \U12/Z_4 ,
         \U12/Z_5 , \U12/Z_6 , \U12/Z_7 , \U12/Z_8 , \U12/Z_9 , \U12/Z_10 ,
         \U12/Z_11 , \U12/Z_12 , \U12/Z_13 , \U12/Z_14 , \U12/Z_15 ,
         \U12/Z_16 , \U12/Z_17 , \U12/Z_18 , \U12/Z_19 , \U12/DATA1_0 ,
         \U12/DATA1_1 , \U12/DATA1_2 , \U12/DATA1_3 , \U12/DATA1_4 ,
         \U12/DATA1_5 , \U12/DATA1_6 , \U12/DATA1_7 , \U12/DATA1_8 ,
         \U12/DATA1_9 , \U12/DATA1_10 , \U12/DATA1_11 , \U12/DATA1_12 ,
         \U12/DATA1_13 , \U12/DATA1_14 , \U12/DATA1_15 , \U12/DATA1_16 ,
         \U12/DATA1_17 , \U12/DATA1_18 , \U12/DATA1_19 , \U11/Z_0 , \U11/Z_1 ,
         \U11/Z_2 , \U11/Z_3 , \U11/Z_4 , \U11/DATA1_0 , \U11/DATA1_1 ,
         \U11/DATA1_2 , \U11/DATA1_3 , \U11/DATA1_4 , \U10/Z_1 , \U10/Z_2 ,
         \U10/Z_3 , \U10/Z_4 , \U10/Z_5 , \U10/Z_6 , \U10/Z_7 , \U10/Z_8 ,
         \U10/Z_9 , \U10/Z_10 , \U10/Z_11 , \U10/Z_12 , \U10/Z_13 , \U10/Z_14 ,
         \U10/Z_15 , \U10/Z_16 , \U10/Z_17 , \U10/Z_18 , \U10/Z_19 ,
         \U10/Z_20 , \U10/Z_21 , \U10/Z_22 , \U10/Z_23 , \U10/Z_24 ,
         \U10/Z_25 , \U10/Z_26 , \U10/Z_27 , \U10/DATA1_1 , \U10/DATA1_2 ,
         \U10/DATA1_3 , \U10/DATA1_4 , \U10/DATA1_5 , \U10/DATA1_6 ,
         \U10/DATA1_7 , \U10/DATA1_8 , \U10/DATA1_9 , \U10/DATA1_10 ,
         \U10/DATA1_11 , \U10/DATA1_12 , \U10/DATA1_13 , \U10/DATA1_14 ,
         \U10/DATA1_15 , \U10/DATA1_16 , \U10/DATA1_17 , \U10/DATA1_18 ,
         \U10/DATA1_19 , \U10/DATA1_20 , \U10/DATA1_21 , \U10/DATA1_22 ,
         \U10/DATA1_23 , \U10/DATA1_24 , \U10/DATA1_25 , \U10/DATA1_26 ,
         \U10/DATA1_27 , \U9/Z_0 , \U9/Z_1 , \U9/Z_2 , \U9/Z_3 , \U9/Z_4 ,
         \U9/Z_5 , \U9/Z_6 , \U9/Z_7 , \U9/Z_8 , \U9/Z_9 , \U9/Z_10 ,
         \U9/Z_11 , \U9/Z_12 , \U9/Z_13 , \U9/Z_14 , \U9/Z_15 , \U9/Z_16 ,
         \U9/Z_17 , \U9/Z_18 , \U9/Z_19 , \U9/DATA1_0 , \U9/DATA1_1 ,
         \U9/DATA1_2 , \U9/DATA1_3 , \U9/DATA1_4 , \U9/DATA1_5 , \U9/DATA1_6 ,
         \U9/DATA1_7 , \U9/DATA1_8 , \U9/DATA1_9 , \U9/DATA1_10 ,
         \U9/DATA1_11 , \U9/DATA1_12 , \U9/DATA1_13 , \U9/DATA1_14 ,
         \U9/DATA1_15 , \U9/DATA1_16 , \U9/DATA1_17 , \U9/DATA1_18 ,
         \U9/DATA1_19 , \U8/Z_0 , \U8/Z_1 , \U8/Z_2 , \U8/Z_3 , \U8/Z_4 ,
         \U8/Z_5 , \U8/DATA1_0 , \U8/DATA1_1 , \U8/DATA1_2 , \U8/DATA1_3 ,
         \U8/DATA1_4 , \U8/DATA1_5 , \U7/Z_1 , \U7/Z_2 , \U7/Z_3 , \U7/Z_4 ,
         \U7/Z_5 , \U7/Z_6 , \U7/Z_7 , \U7/Z_8 , \U7/Z_9 , \U7/Z_10 ,
         \U7/Z_11 , \U7/Z_12 , \U7/Z_13 , \U7/Z_14 , \U7/Z_15 , \U7/Z_16 ,
         \U7/Z_17 , \U7/Z_18 , \U7/Z_19 , \U7/Z_20 , \U7/Z_21 , \U7/Z_22 ,
         \U7/Z_23 , \U7/Z_24 , \U7/Z_25 , \U7/Z_26 , \U7/Z_27 , \U7/DATA1_1 ,
         \U7/DATA1_2 , \U7/DATA1_3 , \U7/DATA1_4 , \U7/DATA1_5 , \U7/DATA1_6 ,
         \U7/DATA1_7 , \U7/DATA1_8 , \U7/DATA1_9 , \U7/DATA1_10 ,
         \U7/DATA1_11 , \U7/DATA1_12 , \U7/DATA1_13 , \U7/DATA1_14 ,
         \U7/DATA1_15 , \U7/DATA1_16 , \U7/DATA1_17 , \U7/DATA1_18 ,
         \U7/DATA1_19 , \U7/DATA1_20 , \U7/DATA1_21 , \U7/DATA1_22 ,
         \U7/DATA1_23 , \U7/DATA1_24 , \U7/DATA1_25 , \U7/DATA1_26 ,
         \U7/DATA1_27 , \U6/Z_0 , \U6/Z_1 , \U6/Z_2 , \U6/Z_3 , \U6/Z_4 ,
         \U6/Z_5 , \U6/Z_6 , \U6/Z_7 , \U6/Z_8 , \U6/Z_9 , \U6/Z_10 ,
         \U6/Z_11 , \U6/Z_12 , \U6/Z_13 , \U6/Z_14 , \U6/Z_15 , \U6/Z_16 ,
         \U6/Z_17 , \U6/Z_18 , \U6/Z_19 , \U6/DATA1_0 , \U6/DATA1_1 ,
         \U6/DATA1_2 , \U6/DATA1_3 , \U6/DATA1_4 , \U6/DATA1_5 , \U6/DATA1_6 ,
         \U6/DATA1_7 , \U6/DATA1_8 , \U6/DATA1_9 , \U6/DATA1_10 ,
         \U6/DATA1_11 , \U6/DATA1_12 , \U6/DATA1_13 , \U6/DATA1_14 ,
         \U6/DATA1_15 , \U6/DATA1_16 , \U6/DATA1_17 , \U6/DATA1_18 ,
         \U6/DATA1_19 , \U5/Z_0 , \U5/Z_1 , \U5/Z_2 , \U5/Z_3 , \U5/Z_4 ,
         \U5/Z_5 , \U5/Z_6 , \U5/DATA1_0 , \U5/DATA1_1 , \U5/DATA1_2 ,
         \U5/DATA1_3 , \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 , \U4/Z_0 ,
         \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 , \U4/Z_7 ,
         \U4/DATA1_0 , \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 , \U4/DATA1_4 ,
         \U4/DATA1_5 , \U4/DATA1_6 , \U4/DATA1_7 , n41, n1092, n1093, n1094,
         n1095, n1096, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;
  assign q[0] = \U4/Z_0 ;
  assign q[1] = \U4/Z_1 ;
  assign q[2] = \U4/Z_2 ;
  assign q[3] = \U4/Z_3 ;
  assign q[4] = \U4/Z_4 ;
  assign q[5] = \U4/Z_5 ;
  assign q[6] = \U4/Z_6 ;
  assign q[7] = \U4/Z_7 ;

  SDFFR_X2 \pipe0_divisor_n_reg[19]  ( .D(1'b0), .SI(n1131), .SE(n1121), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_19 ), .QN(n1118) );
  SDFFR_X2 \pipe0_divisor_n_reg[18]  ( .D(1'b0), .SI(start), .SE(n1127), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_18 ), .QN(n1115) );
  SDFFR_X2 \pipe0_divisor_n_reg[17]  ( .D(1'b0), .SI(start), .SE(n1126), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_17 ), .QN(n1117) );
  SDFFR_X2 \pipe0_divisor_n_reg[16]  ( .D(1'b0), .SI(start), .SE(n1247), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_16 ), .QN(n1116) );
  SDFFR_X2 \pipe0_divisor_n_reg[15]  ( .D(1'b0), .SI(start), .SE(n1248), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_15 ), .QN(n1114) );
  SDFFR_X2 \pipe0_divisor_n_reg[14]  ( .D(1'b0), .SI(n1131), .SE(n1249), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_14 ), .QN(n1113) );
  SDFFR_X2 \pipe0_divisor_n_reg[13]  ( .D(1'b0), .SI(start), .SE(n1123), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_13 ), .QN(n1112) );
  SDFFR_X2 \pipe0_divisor_n_reg[12]  ( .D(1'b0), .SI(start), .SE(n1251), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_12 ), .QN(n1111) );
  SDFFR_X2 \pipe0_divisor_n_reg[11]  ( .D(1'b0), .SI(start), .SE(n1252), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_11 ), .QN(n1110) );
  SDFFR_X2 \pipe0_divisor_n_reg[10]  ( .D(1'b0), .SI(n1131), .SE(n1253), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_10 ), .QN(n1109) );
  SDFFR_X2 \pipe0_divisor_n_reg[9]  ( .D(1'b0), .SI(n1131), .SE(n1120), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_9 ), .QN(n1108) );
  SDFFR_X2 \pipe0_divisor_n_reg[8]  ( .D(1'b0), .SI(n1131), .SE(n1255), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_8 ), .QN(n1107) );
  SDFFR_X2 \pipe0_divisor_n_reg[7]  ( .D(1'b0), .SI(n1131), .SE(n1256), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_7 ), .QN(n1106) );
  SDFFR_X2 \pipe0_divisor_n_reg[6]  ( .D(1'b0), .SI(n1131), .SE(n1257), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_6 ), .QN(n1105) );
  SDFFR_X2 \pipe0_divisor_n_reg[5]  ( .D(1'b0), .SI(n1131), .SE(n1258), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_5 ), .QN(n1104) );
  SDFFR_X2 \pipe0_divisor_n_reg[4]  ( .D(1'b0), .SI(n1131), .SE(n1125), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_4 ), .QN(n1103) );
  SDFFR_X2 \pipe0_divisor_n_reg[3]  ( .D(1'b0), .SI(n1131), .SE(n1260), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_3 ), .QN(n1102) );
  SDFFR_X2 \pipe0_divisor_n_reg[2]  ( .D(1'b0), .SI(n1131), .SE(n1261), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_2 ), .QN(n1101) );
  SDFFR_X2 \pipe0_divisor_n_reg[1]  ( .D(1'b0), .SI(n1131), .SE(n1262), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_1 ), .QN(n1100) );
  SDFFR_X2 \pipe0_divisor_n_reg[0]  ( .D(1'b0), .SI(n1131), .SE(n1263), .CK(
        clock), .RN(n1157), .Q(\U21/DATA1_0 ), .QN(n1099) );
  DFFR_X1 \pipe1_result_reg[27]  ( .D(\U22/Z_27 ), .CK(clock), .RN(n1153), .Q(
        n835) );
  DFFR_X1 \pipe1_result_reg[26]  ( .D(\U22/Z_26 ), .CK(clock), .RN(n1153), .Q(
        n834) );
  DFFR_X1 \pipe1_result_reg[25]  ( .D(\U22/Z_25 ), .CK(clock), .RN(n1153), .Q(
        n833) );
  DFFR_X1 \pipe1_result_reg[24]  ( .D(\U22/Z_24 ), .CK(clock), .RN(n1153), .Q(
        n832) );
  DFFR_X1 \pipe1_result_reg[23]  ( .D(\U22/Z_23 ), .CK(clock), .RN(n1153), .Q(
        n831) );
  DFFR_X1 \pipe1_result_reg[22]  ( .D(\U22/Z_22 ), .CK(clock), .RN(n1153), .Q(
        n830) );
  DFFR_X1 \pipe1_result_reg[21]  ( .D(\U22/Z_21 ), .CK(clock), .RN(n1153), .Q(
        n829) );
  DFFR_X1 \pipe1_result_reg[20]  ( .D(\U22/Z_20 ), .CK(clock), .RN(n1153), .Q(
        n828) );
  DFFR_X1 \pipe1_result_reg[19]  ( .D(\U22/Z_19 ), .CK(clock), .RN(n1153), .Q(
        n827) );
  DFFR_X1 \pipe1_result_reg[17]  ( .D(\U22/Z_17 ), .CK(clock), .RN(n1152), .Q(
        n825) );
  DFFR_X1 \pipe1_result_reg[16]  ( .D(\U22/Z_16 ), .CK(clock), .RN(n1152), .Q(
        n824) );
  DFFR_X1 \pipe1_result_reg[12]  ( .D(\U22/Z_12 ), .CK(clock), .RN(n1152), .Q(
        n820) );
  DFFR_X1 \pipe1_result_reg[11]  ( .D(\U22/Z_11 ), .CK(clock), .RN(n1152), .Q(
        n819) );
  DFFR_X1 \pipe1_result_reg[8]  ( .D(\U22/Z_8 ), .CK(clock), .RN(n1152), .Q(
        n816) );
  DFFR_X1 \pipe1_result_reg[1]  ( .D(\U22/Z_1 ), .CK(clock), .RN(n1151), .Q(
        n809) );
  DFFR_X1 \pipe2_result_reg[27]  ( .D(\U19/Z_27 ), .CK(clock), .RN(n1149), .Q(
        n704) );
  DFFR_X1 \pipe2_result_reg[26]  ( .D(\U19/Z_26 ), .CK(clock), .RN(n1149), .Q(
        n703) );
  DFFR_X1 \pipe2_result_reg[25]  ( .D(\U19/Z_25 ), .CK(clock), .RN(n1149), .Q(
        n702) );
  DFFR_X1 \pipe2_result_reg[24]  ( .D(\U19/Z_24 ), .CK(clock), .RN(n1149), .Q(
        n701) );
  DFFR_X1 \pipe2_result_reg[23]  ( .D(\U19/Z_23 ), .CK(clock), .RN(n1149), .Q(
        n700) );
  DFFR_X1 \pipe2_result_reg[22]  ( .D(\U19/Z_22 ), .CK(clock), .RN(n1149), .Q(
        n699) );
  DFFR_X1 \pipe2_result_reg[21]  ( .D(\U19/Z_21 ), .CK(clock), .RN(n1148), .Q(
        n698) );
  DFFR_X1 \pipe2_result_reg[20]  ( .D(\U19/Z_20 ), .CK(clock), .RN(n1148), .Q(
        n697) );
  DFFR_X1 \pipe2_result_reg[19]  ( .D(\U19/Z_19 ), .CK(clock), .RN(n1148), .Q(
        n696) );
  DFFR_X1 \pipe2_result_reg[18]  ( .D(\U19/Z_18 ), .CK(clock), .RN(n1148), .Q(
        n695) );
  DFFR_X1 \pipe2_result_reg[17]  ( .D(\U19/Z_17 ), .CK(clock), .RN(n1148), .Q(
        n694) );
  DFFR_X1 \pipe2_result_reg[16]  ( .D(\U19/Z_16 ), .CK(clock), .RN(n1148), .Q(
        n693) );
  DFFR_X1 \pipe2_result_reg[15]  ( .D(\U19/Z_15 ), .CK(clock), .RN(n1148), .Q(
        n692) );
  DFFR_X1 \pipe2_result_reg[14]  ( .D(\U19/Z_14 ), .CK(clock), .RN(n1148), .Q(
        n691) );
  DFFR_X1 \pipe2_result_reg[13]  ( .D(\U19/Z_13 ), .CK(clock), .RN(n1148), .Q(
        n690) );
  DFFR_X1 \pipe2_result_reg[12]  ( .D(\U19/Z_12 ), .CK(clock), .RN(n1148), .Q(
        n689) );
  DFFR_X1 \pipe2_result_reg[11]  ( .D(\U19/Z_11 ), .CK(clock), .RN(n1148), .Q(
        n688) );
  DFFR_X1 \pipe2_result_reg[10]  ( .D(\U19/Z_10 ), .CK(clock), .RN(n1148), .Q(
        n687) );
  DFFR_X1 \pipe2_result_reg[9]  ( .D(\U19/Z_9 ), .CK(clock), .RN(n1147), .Q(
        n686) );
  DFFR_X1 \pipe2_result_reg[8]  ( .D(\U19/Z_8 ), .CK(clock), .RN(n1147), .Q(
        n685) );
  DFFR_X1 \pipe2_result_reg[1]  ( .D(\U19/Z_1 ), .CK(clock), .RN(n1147), .Q(
        n678) );
  DFFR_X1 \pipe3_result_reg[27]  ( .D(\U16/Z_27 ), .CK(clock), .RN(n1145), .Q(
        n571) );
  DFFR_X1 \pipe3_result_reg[26]  ( .D(\U16/Z_26 ), .CK(clock), .RN(n1144), .Q(
        n570) );
  DFFR_X1 \pipe3_result_reg[25]  ( .D(\U16/Z_25 ), .CK(clock), .RN(n1144), .Q(
        n569) );
  DFFR_X1 \pipe3_result_reg[24]  ( .D(\U16/Z_24 ), .CK(clock), .RN(n1144), .Q(
        n568) );
  DFFR_X1 \pipe3_result_reg[23]  ( .D(\U16/Z_23 ), .CK(clock), .RN(n1144), .Q(
        n567) );
  DFFR_X1 \pipe3_result_reg[22]  ( .D(\U16/Z_22 ), .CK(clock), .RN(n1144), .Q(
        n566) );
  DFFR_X1 \pipe3_result_reg[21]  ( .D(\U16/Z_21 ), .CK(clock), .RN(n1144), .Q(
        n565) );
  DFFR_X1 \pipe3_result_reg[20]  ( .D(\U16/Z_20 ), .CK(clock), .RN(n1144), .Q(
        n564) );
  DFFR_X1 \pipe3_result_reg[19]  ( .D(\U16/Z_19 ), .CK(clock), .RN(n1144), .Q(
        n563) );
  DFFR_X1 \pipe3_result_reg[18]  ( .D(\U16/Z_18 ), .CK(clock), .RN(n1144), .Q(
        n562) );
  DFFR_X1 \pipe3_result_reg[17]  ( .D(\U16/Z_17 ), .CK(clock), .RN(n1144), .Q(
        n561) );
  DFFR_X1 \pipe3_result_reg[16]  ( .D(\U16/Z_16 ), .CK(clock), .RN(n1144), .Q(
        n560) );
  DFFR_X1 \pipe3_result_reg[15]  ( .D(\U16/Z_15 ), .CK(clock), .RN(n1144), .Q(
        n559) );
  DFFR_X1 \pipe3_result_reg[14]  ( .D(\U16/Z_14 ), .CK(clock), .RN(n1143), .Q(
        n558) );
  DFFR_X1 \pipe3_result_reg[13]  ( .D(\U16/Z_13 ), .CK(clock), .RN(n1143), .Q(
        n557) );
  DFFR_X1 \pipe3_result_reg[12]  ( .D(\U16/Z_12 ), .CK(clock), .RN(n1143), .Q(
        n556) );
  DFFR_X1 \pipe3_result_reg[11]  ( .D(\U16/Z_11 ), .CK(clock), .RN(n1143), .Q(
        n555) );
  DFFR_X1 \pipe3_result_reg[10]  ( .D(\U16/Z_10 ), .CK(clock), .RN(n1143), .Q(
        n554) );
  DFFR_X1 \pipe3_result_reg[9]  ( .D(\U16/Z_9 ), .CK(clock), .RN(n1143), .Q(
        n553) );
  DFFR_X1 \pipe3_result_reg[8]  ( .D(\U16/Z_8 ), .CK(clock), .RN(n1143), .Q(
        n552) );
  DFFR_X1 \pipe3_result_reg[1]  ( .D(\U16/Z_1 ), .CK(clock), .RN(n1142), .Q(
        n545) );
  DFFR_X1 \pipe4_result_reg[27]  ( .D(\U13/Z_27 ), .CK(clock), .RN(n1155), .Q(
        n436) );
  DFFR_X1 \pipe4_result_reg[26]  ( .D(\U13/Z_26 ), .CK(clock), .RN(n1157), .Q(
        n435) );
  DFFR_X1 \pipe4_result_reg[25]  ( .D(\U13/Z_25 ), .CK(clock), .RN(n1156), .Q(
        n434) );
  DFFR_X1 \pipe4_result_reg[24]  ( .D(\U13/Z_24 ), .CK(clock), .RN(n1155), .Q(
        n433) );
  DFFR_X1 \pipe4_result_reg[23]  ( .D(\U13/Z_23 ), .CK(clock), .RN(n1145), .Q(
        n432) );
  DFFR_X1 \pipe4_result_reg[22]  ( .D(\U13/Z_22 ), .CK(clock), .RN(n1156), .Q(
        n431) );
  DFFR_X1 \pipe4_result_reg[21]  ( .D(\U13/Z_21 ), .CK(clock), .RN(n1136), .Q(
        n430) );
  DFFR_X1 \pipe4_result_reg[20]  ( .D(\U13/Z_20 ), .CK(clock), .RN(n1157), .Q(
        n429) );
  DFFR_X1 \pipe4_result_reg[19]  ( .D(\U13/Z_19 ), .CK(clock), .RN(n1134), .Q(
        n428) );
  DFFR_X1 \pipe4_result_reg[18]  ( .D(\U13/Z_18 ), .CK(clock), .RN(reset_n), 
        .Q(n427) );
  DFFR_X1 \pipe4_result_reg[17]  ( .D(\U13/Z_17 ), .CK(clock), .RN(n1143), .Q(
        n426) );
  DFFR_X1 \pipe4_result_reg[16]  ( .D(\U13/Z_16 ), .CK(clock), .RN(n1139), .Q(
        n425) );
  DFFR_X1 \pipe4_result_reg[15]  ( .D(\U13/Z_15 ), .CK(clock), .RN(n1149), .Q(
        n424) );
  DFFR_X1 \pipe4_result_reg[14]  ( .D(\U13/Z_14 ), .CK(clock), .RN(n1144), .Q(
        n423) );
  DFFR_X1 \pipe4_result_reg[13]  ( .D(\U13/Z_13 ), .CK(clock), .RN(n1148), .Q(
        n422) );
  DFFR_X1 \pipe4_result_reg[12]  ( .D(\U13/Z_12 ), .CK(clock), .RN(n1152), .Q(
        n421) );
  DFFR_X1 \pipe4_result_reg[11]  ( .D(\U13/Z_11 ), .CK(clock), .RN(n1135), .Q(
        n420) );
  DFFR_X1 \pipe4_result_reg[10]  ( .D(\U13/Z_10 ), .CK(clock), .RN(n1153), .Q(
        n419) );
  DFFR_X1 \pipe4_result_reg[9]  ( .D(\U13/Z_9 ), .CK(clock), .RN(n1138), .Q(
        n418) );
  DFFR_X1 \pipe4_result_reg[8]  ( .D(\U13/Z_8 ), .CK(clock), .RN(n1141), .Q(
        n417) );
  DFFR_X1 \pipe4_result_reg[1]  ( .D(\U13/Z_1 ), .CK(clock), .RN(n1141), .Q(
        n410) );
  DFFR_X1 \pipe5_result_reg[27]  ( .D(\U10/Z_27 ), .CK(clock), .RN(n1139), .Q(
        n299) );
  DFFR_X1 \pipe5_result_reg[26]  ( .D(\U10/Z_26 ), .CK(clock), .RN(n1139), .Q(
        n298) );
  DFFR_X1 \pipe5_result_reg[25]  ( .D(\U10/Z_25 ), .CK(clock), .RN(n1139), .Q(
        n297) );
  DFFR_X1 \pipe5_result_reg[24]  ( .D(\U10/Z_24 ), .CK(clock), .RN(n1139), .Q(
        n296) );
  DFFR_X1 \pipe5_result_reg[23]  ( .D(\U10/Z_23 ), .CK(clock), .RN(n1139), .Q(
        n295) );
  DFFR_X1 \pipe5_result_reg[22]  ( .D(\U10/Z_22 ), .CK(clock), .RN(n1139), .Q(
        n294) );
  DFFR_X1 \pipe5_result_reg[21]  ( .D(\U10/Z_21 ), .CK(clock), .RN(n1139), .Q(
        n293) );
  DFFR_X1 \pipe5_result_reg[20]  ( .D(\U10/Z_20 ), .CK(clock), .RN(n1139), .Q(
        n292) );
  DFFR_X1 \pipe5_result_reg[19]  ( .D(\U10/Z_19 ), .CK(clock), .RN(n1139), .Q(
        n291) );
  DFFR_X1 \pipe5_result_reg[18]  ( .D(\U10/Z_18 ), .CK(clock), .RN(n1139), .Q(
        n290) );
  DFFR_X1 \pipe5_result_reg[17]  ( .D(\U10/Z_17 ), .CK(clock), .RN(n1139), .Q(
        n289) );
  DFFR_X1 \pipe5_result_reg[16]  ( .D(\U10/Z_16 ), .CK(clock), .RN(n1139), .Q(
        n288) );
  DFFR_X1 \pipe5_result_reg[15]  ( .D(\U10/Z_15 ), .CK(clock), .RN(n1138), .Q(
        n287) );
  DFFR_X1 \pipe5_result_reg[14]  ( .D(\U10/Z_14 ), .CK(clock), .RN(n1138), .Q(
        n286) );
  DFFR_X1 \pipe5_result_reg[13]  ( .D(\U10/Z_13 ), .CK(clock), .RN(n1138), .Q(
        n285) );
  DFFR_X1 \pipe5_result_reg[12]  ( .D(\U10/Z_12 ), .CK(clock), .RN(n1138), .Q(
        n284) );
  DFFR_X1 \pipe5_result_reg[11]  ( .D(\U10/Z_11 ), .CK(clock), .RN(n1138), .Q(
        n283) );
  DFFR_X1 \pipe5_result_reg[10]  ( .D(\U10/Z_10 ), .CK(clock), .RN(n1138), .Q(
        n282) );
  DFFR_X1 \pipe5_result_reg[9]  ( .D(\U10/Z_9 ), .CK(clock), .RN(n1138), .Q(
        n281) );
  DFFR_X1 \pipe5_result_reg[8]  ( .D(\U10/Z_8 ), .CK(clock), .RN(n1138), .Q(
        n280) );
  DFFR_X1 \pipe5_result_reg[1]  ( .D(\U10/Z_1 ), .CK(clock), .RN(n1137), .Q(
        n273) );
  DFFR_X1 \pipe6_result_reg[27]  ( .D(\U7/Z_27 ), .CK(clock), .RN(n1135), .Q(
        n160) );
  DFFR_X1 \pipe6_result_reg[26]  ( .D(\U7/Z_26 ), .CK(clock), .RN(n1135), .Q(
        n159) );
  DFFR_X1 \pipe6_result_reg[25]  ( .D(\U7/Z_25 ), .CK(clock), .RN(n1135), .Q(
        n158) );
  DFFR_X1 \pipe6_result_reg[24]  ( .D(\U7/Z_24 ), .CK(clock), .RN(n1135), .Q(
        n157) );
  DFFR_X1 \pipe6_result_reg[23]  ( .D(\U7/Z_23 ), .CK(clock), .RN(n1134), .Q(
        n156) );
  DFFR_X1 \pipe6_result_reg[22]  ( .D(\U7/Z_22 ), .CK(clock), .RN(n1134), .Q(
        n155) );
  DFFR_X1 \pipe6_result_reg[21]  ( .D(\U7/Z_21 ), .CK(clock), .RN(n1134), .Q(
        n154) );
  DFFR_X1 \pipe6_result_reg[20]  ( .D(\U7/Z_20 ), .CK(clock), .RN(n1134), .Q(
        n153) );
  DFFR_X1 \pipe6_result_reg[19]  ( .D(\U7/Z_19 ), .CK(clock), .RN(n1134), .Q(
        n152) );
  DFFR_X1 \pipe6_result_reg[18]  ( .D(\U7/Z_18 ), .CK(clock), .RN(n1134), .Q(
        n151) );
  DFFR_X1 \pipe6_result_reg[17]  ( .D(\U7/Z_17 ), .CK(clock), .RN(n1134), .Q(
        n150) );
  DFFR_X1 \pipe6_result_reg[16]  ( .D(\U7/Z_16 ), .CK(clock), .RN(n1134), .Q(
        n149) );
  DFFR_X1 \pipe6_result_reg[15]  ( .D(\U7/Z_15 ), .CK(clock), .RN(n1134), .Q(
        n148) );
  DFFR_X1 \pipe6_result_reg[14]  ( .D(\U7/Z_14 ), .CK(clock), .RN(n1134), .Q(
        n147) );
  DFFR_X1 \pipe6_result_reg[13]  ( .D(\U7/Z_13 ), .CK(clock), .RN(n1134), .Q(
        n146) );
  DFFR_X1 \pipe6_result_reg[12]  ( .D(\U7/Z_12 ), .CK(clock), .RN(n1134), .Q(
        n145) );
  DFFR_X1 \pipe6_result_reg[10]  ( .D(\U7/Z_10 ), .CK(clock), .RN(n1133), .Q(
        n143) );
  DFFR_X1 \pipe6_result_reg[9]  ( .D(\U7/Z_9 ), .CK(clock), .RN(n1133), .Q(
        n142) );
  DFFR_X1 \pipe6_result_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .RN(n1133), .Q(
        n134) );
  AND2_X1 U56 ( .A1(\U9/DATA1_19 ), .A2(n383), .ZN(\U9/Z_19 ) );
  AND2_X1 U57 ( .A1(\U9/DATA1_18 ), .A2(n383), .ZN(\U9/Z_18 ) );
  AND2_X1 U58 ( .A1(\U9/DATA1_17 ), .A2(n383), .ZN(\U9/Z_17 ) );
  AND2_X1 U59 ( .A1(\U9/DATA1_16 ), .A2(n383), .ZN(\U9/Z_16 ) );
  AND2_X1 U68 ( .A1(\U8/DATA1_5 ), .A2(n383), .ZN(\U8/Z_5 ) );
  AND2_X1 U69 ( .A1(\U8/DATA1_4 ), .A2(n383), .ZN(\U8/Z_4 ) );
  AND2_X1 U70 ( .A1(\U8/DATA1_3 ), .A2(n383), .ZN(\U8/Z_3 ) );
  AND2_X1 U71 ( .A1(\U8/DATA1_2 ), .A2(n383), .ZN(\U8/Z_2 ) );
  AND2_X1 U77 ( .A1(\U7/DATA1_6 ), .A2(n245), .ZN(\U7/Z_6 ) );
  AND2_X1 U78 ( .A1(\U7/DATA1_5 ), .A2(n245), .ZN(\U7/Z_5 ) );
  AND2_X1 U79 ( .A1(\U7/DATA1_4 ), .A2(n245), .ZN(\U7/Z_4 ) );
  AND2_X1 U80 ( .A1(\U7/DATA1_3 ), .A2(n245), .ZN(\U7/Z_3 ) );
  AND2_X1 U89 ( .A1(\U7/DATA1_2 ), .A2(n245), .ZN(\U7/Z_2 ) );
  AND2_X1 U100 ( .A1(\U7/DATA1_1 ), .A2(n245), .ZN(\U7/Z_1 ) );
  AND2_X1 U110 ( .A1(\U6/DATA1_19 ), .A2(n245), .ZN(\U6/Z_19 ) );
  AND2_X1 U111 ( .A1(\U6/DATA1_18 ), .A2(n245), .ZN(\U6/Z_18 ) );
  AND2_X1 U112 ( .A1(\U6/DATA1_17 ), .A2(n245), .ZN(\U6/Z_17 ) );
  AND2_X1 U113 ( .A1(\U6/DATA1_16 ), .A2(n245), .ZN(\U6/Z_16 ) );
  AND2_X1 U122 ( .A1(\U5/DATA1_6 ), .A2(n245), .ZN(\U5/Z_6 ) );
  AND2_X1 U123 ( .A1(\U5/DATA1_5 ), .A2(n245), .ZN(\U5/Z_5 ) );
  AND2_X1 U124 ( .A1(\U5/DATA1_4 ), .A2(n245), .ZN(\U5/Z_4 ) );
  AND2_X1 U125 ( .A1(\U5/DATA1_3 ), .A2(n245), .ZN(\U5/Z_3 ) );
  AND2_X1 U126 ( .A1(\U5/DATA1_2 ), .A2(n245), .ZN(\U5/Z_2 ) );
  AND2_X1 U129 ( .A1(\U4/DATA1_7 ), .A2(n41), .ZN(\U4/Z_7 ) );
  AND2_X1 U130 ( .A1(\U4/DATA1_6 ), .A2(n41), .ZN(\U4/Z_6 ) );
  AND2_X1 U131 ( .A1(\U4/DATA1_5 ), .A2(n41), .ZN(\U4/Z_5 ) );
  AND2_X1 U132 ( .A1(\U4/DATA1_4 ), .A2(n41), .ZN(\U4/Z_4 ) );
  AND2_X1 U133 ( .A1(\U4/DATA1_3 ), .A2(n41), .ZN(\U4/Z_3 ) );
  AND2_X1 U134 ( .A1(\U4/DATA1_2 ), .A2(n41), .ZN(\U4/Z_2 ) );
  AND2_X1 U144 ( .A1(\U25/DATA1_6 ), .A2(start), .ZN(\U25/Z_6 ) );
  AND2_X1 U145 ( .A1(\U25/DATA1_5 ), .A2(start), .ZN(\U25/Z_5 ) );
  AND2_X1 U146 ( .A1(\U25/DATA1_4 ), .A2(start), .ZN(\U25/Z_4 ) );
  AND2_X1 U147 ( .A1(\U25/DATA1_3 ), .A2(start), .ZN(\U25/Z_3 ) );
  AND2_X1 U156 ( .A1(\U25/DATA1_2 ), .A2(start), .ZN(\U25/Z_2 ) );
  AND2_X1 U167 ( .A1(\U25/DATA1_1 ), .A2(n1131), .ZN(\U25/Z_1 ) );
  AND2_X1 U173 ( .A1(\U22/DATA1_6 ), .A2(n915), .ZN(\U22/Z_6 ) );
  AND2_X1 U174 ( .A1(\U22/DATA1_5 ), .A2(n915), .ZN(\U22/Z_5 ) );
  AND2_X1 U175 ( .A1(\U22/DATA1_4 ), .A2(n915), .ZN(\U22/Z_4 ) );
  AND2_X1 U176 ( .A1(\U22/DATA1_3 ), .A2(n915), .ZN(\U22/Z_3 ) );
  AND2_X1 U185 ( .A1(\U22/DATA1_2 ), .A2(n915), .ZN(\U22/Z_2 ) );
  AND2_X1 U196 ( .A1(\U22/DATA1_1 ), .A2(n915), .ZN(\U22/Z_1 ) );
  AND2_X1 U223 ( .A1(\U19/DATA1_6 ), .A2(n1098), .ZN(\U19/Z_6 ) );
  AND2_X1 U224 ( .A1(\U19/DATA1_5 ), .A2(n1098), .ZN(\U19/Z_5 ) );
  AND2_X1 U225 ( .A1(\U19/DATA1_4 ), .A2(n1098), .ZN(\U19/Z_4 ) );
  AND2_X1 U226 ( .A1(\U19/DATA1_3 ), .A2(n1098), .ZN(\U19/Z_3 ) );
  AND2_X1 U235 ( .A1(\U19/DATA1_2 ), .A2(n1098), .ZN(\U19/Z_2 ) );
  AND2_X1 U246 ( .A1(\U19/DATA1_1 ), .A2(n1098), .ZN(\U19/Z_1 ) );
  AND2_X1 U256 ( .A1(\U18/DATA1_19 ), .A2(n1098), .ZN(\U18/Z_19 ) );
  AND2_X1 U257 ( .A1(\U18/DATA1_18 ), .A2(n1098), .ZN(\U18/Z_18 ) );
  AND2_X1 U258 ( .A1(\U18/DATA1_17 ), .A2(n1098), .ZN(\U18/Z_17 ) );
  AND2_X1 U259 ( .A1(\U18/DATA1_16 ), .A2(n1098), .ZN(\U18/Z_16 ) );
  AND2_X1 U268 ( .A1(\U17/DATA1_2 ), .A2(n1098), .ZN(\U17/Z_2 ) );
  AND2_X1 U274 ( .A1(\U16/DATA1_6 ), .A2(n653), .ZN(\U16/Z_6 ) );
  AND2_X1 U275 ( .A1(\U16/DATA1_5 ), .A2(n653), .ZN(\U16/Z_5 ) );
  AND2_X1 U276 ( .A1(\U16/DATA1_4 ), .A2(n653), .ZN(\U16/Z_4 ) );
  AND2_X1 U277 ( .A1(\U16/DATA1_3 ), .A2(n653), .ZN(\U16/Z_3 ) );
  AND2_X1 U286 ( .A1(\U16/DATA1_2 ), .A2(n653), .ZN(\U16/Z_2 ) );
  AND2_X1 U297 ( .A1(\U16/DATA1_1 ), .A2(n653), .ZN(\U16/Z_1 ) );
  AND2_X1 U307 ( .A1(\U15/DATA1_19 ), .A2(n653), .ZN(\U15/Z_19 ) );
  AND2_X1 U308 ( .A1(\U15/DATA1_18 ), .A2(n653), .ZN(\U15/Z_18 ) );
  AND2_X1 U309 ( .A1(\U15/DATA1_17 ), .A2(n653), .ZN(\U15/Z_17 ) );
  AND2_X1 U310 ( .A1(\U15/DATA1_16 ), .A2(n653), .ZN(\U15/Z_16 ) );
  AND2_X1 U319 ( .A1(\U14/DATA1_3 ), .A2(n653), .ZN(\U14/Z_3 ) );
  AND2_X1 U320 ( .A1(\U14/DATA1_2 ), .A2(n653), .ZN(\U14/Z_2 ) );
  AND2_X1 U326 ( .A1(\U13/DATA1_6 ), .A2(n519), .ZN(\U13/Z_6 ) );
  AND2_X1 U327 ( .A1(\U13/DATA1_5 ), .A2(n519), .ZN(\U13/Z_5 ) );
  AND2_X1 U328 ( .A1(\U13/DATA1_4 ), .A2(n519), .ZN(\U13/Z_4 ) );
  AND2_X1 U329 ( .A1(\U13/DATA1_3 ), .A2(n519), .ZN(\U13/Z_3 ) );
  AND2_X1 U338 ( .A1(\U13/DATA1_2 ), .A2(n519), .ZN(\U13/Z_2 ) );
  AND2_X1 U349 ( .A1(\U13/DATA1_1 ), .A2(n519), .ZN(\U13/Z_1 ) );
  AND2_X1 U359 ( .A1(\U12/DATA1_19 ), .A2(n519), .ZN(\U12/Z_19 ) );
  AND2_X1 U360 ( .A1(\U12/DATA1_18 ), .A2(n519), .ZN(\U12/Z_18 ) );
  AND2_X1 U361 ( .A1(\U12/DATA1_17 ), .A2(n519), .ZN(\U12/Z_17 ) );
  AND2_X1 U362 ( .A1(\U12/DATA1_16 ), .A2(n519), .ZN(\U12/Z_16 ) );
  AND2_X1 U371 ( .A1(\U11/DATA1_4 ), .A2(n519), .ZN(\U11/Z_4 ) );
  AND2_X1 U372 ( .A1(\U11/DATA1_3 ), .A2(n519), .ZN(\U11/Z_3 ) );
  AND2_X1 U373 ( .A1(\U11/DATA1_2 ), .A2(n519), .ZN(\U11/Z_2 ) );
  AND2_X1 U379 ( .A1(\U10/DATA1_6 ), .A2(n383), .ZN(\U10/Z_6 ) );
  AND2_X1 U380 ( .A1(\U10/DATA1_5 ), .A2(n383), .ZN(\U10/Z_5 ) );
  AND2_X1 U381 ( .A1(\U10/DATA1_4 ), .A2(n383), .ZN(\U10/Z_4 ) );
  AND2_X1 U382 ( .A1(\U10/DATA1_3 ), .A2(n383), .ZN(\U10/Z_3 ) );
  AND2_X1 U391 ( .A1(\U10/DATA1_2 ), .A2(n383), .ZN(\U10/Z_2 ) );
  AND2_X1 U402 ( .A1(\U10/DATA1_1 ), .A2(n383), .ZN(\U10/Z_1 ) );
  pipleline_stage_1 stage0 ( .divided(divided), .divisor({n1121, n1127, n1126, 
        n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
        n1257, n1258, n1259, n1260, n1261, n1262, n1263}), .q(\U23/DATA1_0 ), 
        .stage_out({\U25/DATA1_27 , \U25/DATA1_26 , \U25/DATA1_25 , 
        \U25/DATA1_24 , \U25/DATA1_23 , \U25/DATA1_22 , \U25/DATA1_21 , 
        \U25/DATA1_20 , \U25/DATA1_19 , \U25/DATA1_18 , \U25/DATA1_17 , 
        \U25/DATA1_16 , \U25/DATA1_15 , \U25/DATA1_14 , \U25/DATA1_13 , 
        \U25/DATA1_12 , \U25/DATA1_11 , \U25/DATA1_10 , \U25/DATA1_9 , 
        \U25/DATA1_8 , \U25/DATA1_7 , \U25/DATA1_6 , \U25/DATA1_5 , 
        \U25/DATA1_4 , \U25/DATA1_3 , \U25/DATA1_2 , \U25/DATA1_1 , 
        SYNOPSYS_UNCONNECTED__0}) );
  pipleline_stage_7 stage1 ( .divided({n964, n963, n962, n961, n960, n959, 
        n958, n957, n956, n955, n954, n953, n952, n951, n950, n949, n948, n947, 
        n946, n945, n944, n943, n942, n941, n940, n939, n938, 1'b0}), 
        .divisor({\U21/DATA1_19 , \U21/DATA1_18 , \U21/DATA1_17 , 
        \U21/DATA1_16 , \U21/DATA1_15 , \U21/DATA1_14 , \U21/DATA1_13 , 
        \U21/DATA1_12 , \U21/DATA1_11 , \U21/DATA1_10 , \U21/DATA1_9 , 
        \U21/DATA1_8 , \U21/DATA1_7 , \U21/DATA1_6 , \U21/DATA1_5 , 
        \U21/DATA1_4 , \U21/DATA1_3 , \U21/DATA1_2 , \U21/DATA1_1 , 
        \U21/DATA1_0 }), .q(\U20/DATA1_0 ), .stage_out({\U22/DATA1_27 , 
        \U22/DATA1_26 , \U22/DATA1_25 , \U22/DATA1_24 , \U22/DATA1_23 , 
        \U22/DATA1_22 , \U22/DATA1_21 , \U22/DATA1_20 , \U22/DATA1_19 , 
        \U22/DATA1_18 , \U22/DATA1_17 , \U22/DATA1_16 , \U22/DATA1_15 , 
        \U22/DATA1_14 , \U22/DATA1_13 , \U22/DATA1_12 , \U22/DATA1_11 , 
        \U22/DATA1_10 , \U22/DATA1_9 , \U22/DATA1_8 , \U22/DATA1_7 , 
        \U22/DATA1_6 , \U22/DATA1_5 , \U22/DATA1_4 , \U22/DATA1_3 , 
        \U22/DATA1_2 , \U22/DATA1_1 , SYNOPSYS_UNCONNECTED__1}) );
  pipleline_stage_6 stage2 ( .divided({n835, n834, n833, n832, n831, n830, 
        n829, n828, n827, n826, n825, n824, n823, n822, n821, n820, n819, n818, 
        n817, n816, n815, n814, n813, n812, n811, n810, n809, 1'b0}), 
        .divisor({\U18/DATA1_19 , \U18/DATA1_18 , \U18/DATA1_17 , 
        \U18/DATA1_16 , \U18/DATA1_15 , \U18/DATA1_14 , \U18/DATA1_13 , 
        \U18/DATA1_12 , \U18/DATA1_11 , \U18/DATA1_10 , \U18/DATA1_9 , 
        \U18/DATA1_8 , \U18/DATA1_7 , \U18/DATA1_6 , \U18/DATA1_5 , 
        \U18/DATA1_4 , \U18/DATA1_3 , \U18/DATA1_2 , \U18/DATA1_1 , 
        \U18/DATA1_0 }), .q(\U17/DATA1_0 ), .stage_out({\U19/DATA1_27 , 
        \U19/DATA1_26 , \U19/DATA1_25 , \U19/DATA1_24 , \U19/DATA1_23 , 
        \U19/DATA1_22 , \U19/DATA1_21 , \U19/DATA1_20 , \U19/DATA1_19 , 
        \U19/DATA1_18 , \U19/DATA1_17 , \U19/DATA1_16 , \U19/DATA1_15 , 
        \U19/DATA1_14 , \U19/DATA1_13 , \U19/DATA1_12 , \U19/DATA1_11 , 
        \U19/DATA1_10 , \U19/DATA1_9 , \U19/DATA1_8 , \U19/DATA1_7 , 
        \U19/DATA1_6 , \U19/DATA1_5 , \U19/DATA1_4 , \U19/DATA1_3 , 
        \U19/DATA1_2 , \U19/DATA1_1 , SYNOPSYS_UNCONNECTED__2}) );
  pipleline_stage_5 stage3 ( .divided({n704, n703, n702, n701, n700, n699, 
        n698, n697, n696, n695, n694, n693, n692, n691, n690, n689, n688, n687, 
        n686, n685, n684, n683, n682, n681, n680, n679, n678, 1'b0}), 
        .divisor({\U15/DATA1_19 , \U15/DATA1_18 , \U15/DATA1_17 , 
        \U15/DATA1_16 , \U15/DATA1_15 , \U15/DATA1_14 , \U15/DATA1_13 , 
        \U15/DATA1_12 , \U15/DATA1_11 , \U15/DATA1_10 , \U15/DATA1_9 , 
        \U15/DATA1_8 , \U15/DATA1_7 , \U15/DATA1_6 , \U15/DATA1_5 , 
        \U15/DATA1_4 , \U15/DATA1_3 , \U15/DATA1_2 , \U15/DATA1_1 , 
        \U15/DATA1_0 }), .q(\U14/DATA1_0 ), .stage_out({\U16/DATA1_27 , 
        \U16/DATA1_26 , \U16/DATA1_25 , \U16/DATA1_24 , \U16/DATA1_23 , 
        \U16/DATA1_22 , \U16/DATA1_21 , \U16/DATA1_20 , \U16/DATA1_19 , 
        \U16/DATA1_18 , \U16/DATA1_17 , \U16/DATA1_16 , \U16/DATA1_15 , 
        \U16/DATA1_14 , \U16/DATA1_13 , \U16/DATA1_12 , \U16/DATA1_11 , 
        \U16/DATA1_10 , \U16/DATA1_9 , \U16/DATA1_8 , \U16/DATA1_7 , 
        \U16/DATA1_6 , \U16/DATA1_5 , \U16/DATA1_4 , \U16/DATA1_3 , 
        \U16/DATA1_2 , \U16/DATA1_1 , SYNOPSYS_UNCONNECTED__3}) );
  pipleline_stage_4 stage4 ( .divided({n571, n570, n569, n568, n567, n566, 
        n565, n564, n563, n562, n561, n560, n559, n558, n557, n556, n555, n554, 
        n553, n552, n551, n550, n549, n548, n547, n546, n545, 1'b0}), 
        .divisor({\U12/DATA1_19 , \U12/DATA1_18 , \U12/DATA1_17 , 
        \U12/DATA1_16 , \U12/DATA1_15 , \U12/DATA1_14 , \U12/DATA1_13 , 
        \U12/DATA1_12 , \U12/DATA1_11 , \U12/DATA1_10 , \U12/DATA1_9 , 
        \U12/DATA1_8 , \U12/DATA1_7 , \U12/DATA1_6 , \U12/DATA1_5 , 
        \U12/DATA1_4 , \U12/DATA1_3 , \U12/DATA1_2 , \U12/DATA1_1 , 
        \U12/DATA1_0 }), .q(\U11/DATA1_0 ), .stage_out({\U13/DATA1_27 , 
        \U13/DATA1_26 , \U13/DATA1_25 , \U13/DATA1_24 , \U13/DATA1_23 , 
        \U13/DATA1_22 , \U13/DATA1_21 , \U13/DATA1_20 , \U13/DATA1_19 , 
        \U13/DATA1_18 , \U13/DATA1_17 , \U13/DATA1_16 , \U13/DATA1_15 , 
        \U13/DATA1_14 , \U13/DATA1_13 , \U13/DATA1_12 , \U13/DATA1_11 , 
        \U13/DATA1_10 , \U13/DATA1_9 , \U13/DATA1_8 , \U13/DATA1_7 , 
        \U13/DATA1_6 , \U13/DATA1_5 , \U13/DATA1_4 , \U13/DATA1_3 , 
        \U13/DATA1_2 , \U13/DATA1_1 , SYNOPSYS_UNCONNECTED__4}) );
  pipleline_stage_3 stage5 ( .divided({n436, n435, n434, n433, n432, n431, 
        n430, n429, n428, n427, n426, n425, n424, n423, n422, n421, n420, n419, 
        n418, n417, n416, n415, n414, n413, n412, n411, n410, 1'b0}), 
        .divisor({\U9/DATA1_19 , \U9/DATA1_18 , \U9/DATA1_17 , \U9/DATA1_16 , 
        \U9/DATA1_15 , \U9/DATA1_14 , \U9/DATA1_13 , \U9/DATA1_12 , 
        \U9/DATA1_11 , \U9/DATA1_10 , \U9/DATA1_9 , \U9/DATA1_8 , \U9/DATA1_7 , 
        \U9/DATA1_6 , \U9/DATA1_5 , \U9/DATA1_4 , \U9/DATA1_3 , \U9/DATA1_2 , 
        \U9/DATA1_1 , \U9/DATA1_0 }), .q(\U8/DATA1_0 ), .stage_out({
        \U10/DATA1_27 , \U10/DATA1_26 , \U10/DATA1_25 , \U10/DATA1_24 , 
        \U10/DATA1_23 , \U10/DATA1_22 , \U10/DATA1_21 , \U10/DATA1_20 , 
        \U10/DATA1_19 , \U10/DATA1_18 , \U10/DATA1_17 , \U10/DATA1_16 , 
        \U10/DATA1_15 , \U10/DATA1_14 , \U10/DATA1_13 , \U10/DATA1_12 , 
        \U10/DATA1_11 , \U10/DATA1_10 , \U10/DATA1_9 , \U10/DATA1_8 , 
        \U10/DATA1_7 , \U10/DATA1_6 , \U10/DATA1_5 , \U10/DATA1_4 , 
        \U10/DATA1_3 , \U10/DATA1_2 , \U10/DATA1_1 , SYNOPSYS_UNCONNECTED__5})
         );
  pipleline_stage_2 stage6 ( .divided({n299, n298, n297, n296, n295, n294, 
        n293, n292, n291, n290, n289, n288, n287, n286, n285, n284, n283, n282, 
        n281, n280, n279, n278, n277, n276, n275, n274, n273, 1'b0}), 
        .divisor({\U6/DATA1_19 , \U6/DATA1_18 , \U6/DATA1_17 , \U6/DATA1_16 , 
        \U6/DATA1_15 , \U6/DATA1_14 , \U6/DATA1_13 , \U6/DATA1_12 , 
        \U6/DATA1_11 , \U6/DATA1_10 , \U6/DATA1_9 , \U6/DATA1_8 , \U6/DATA1_7 , 
        \U6/DATA1_6 , \U6/DATA1_5 , \U6/DATA1_4 , \U6/DATA1_3 , \U6/DATA1_2 , 
        \U6/DATA1_1 , \U6/DATA1_0 }), .q(\U5/DATA1_0 ), .stage_out({
        \U7/DATA1_27 , \U7/DATA1_26 , \U7/DATA1_25 , \U7/DATA1_24 , 
        \U7/DATA1_23 , \U7/DATA1_22 , \U7/DATA1_21 , \U7/DATA1_20 , 
        \U7/DATA1_19 , \U7/DATA1_18 , \U7/DATA1_17 , \U7/DATA1_16 , 
        \U7/DATA1_15 , \U7/DATA1_14 , \U7/DATA1_13 , \U7/DATA1_12 , 
        \U7/DATA1_11 , \U7/DATA1_10 , \U7/DATA1_9 , \U7/DATA1_8 , \U7/DATA1_7 , 
        \U7/DATA1_6 , \U7/DATA1_5 , \U7/DATA1_4 , \U7/DATA1_3 , \U7/DATA1_2 , 
        \U7/DATA1_1 , SYNOPSYS_UNCONNECTED__6}) );
  pipleline_stage_0 stage7 ( .divided({n160, n159, n158, n157, n156, n155, 
        n154, n153, n152, n151, n150, n149, n148, n147, n146, n145, n144, n143, 
        n142, n141, n140, n139, n138, n137, n136, n135, n134, 1'b0}), 
        .divisor({n132, n131, n130, n129, n128, n127, n126, n125, n124, n123, 
        n122, n121, n120, n119, n118, n117, n116, n115, n114, n113}), .q(
        \U4/DATA1_0 ) );
  DFFR_X2 \pipe6_divisor_n_reg[0]  ( .D(\U6/Z_0 ), .CK(clock), .RN(n1136), .Q(
        n113) );
  DFFR_X2 \pipe0_result_reg[20]  ( .D(\U25/Z_20 ), .CK(clock), .RN(n1156), .Q(
        n957) );
  DFFR_X2 \pipe0_result_reg[21]  ( .D(\U25/Z_21 ), .CK(clock), .RN(n1156), .Q(
        n958) );
  DFFR_X2 StartOut1_reg ( .D(n915), .CK(clock), .RN(n1153), .Q(n1098), .QN(
        n1096) );
  DFFR_X2 StartOut0_reg ( .D(start), .CK(clock), .RN(n1157), .Q(n915), .QN(
        n1130) );
  DFFR_X2 \pipe6_divisor_n_reg[15]  ( .D(\U6/Z_15 ), .CK(clock), .RN(n1137), 
        .Q(n128) );
  DFFR_X2 \pipe6_divisor_n_reg[14]  ( .D(\U6/Z_14 ), .CK(clock), .RN(n1137), 
        .Q(n127) );
  DFFR_X2 \pipe5_divisor_n_reg[15]  ( .D(\U9/Z_15 ), .CK(clock), .RN(n1140), 
        .Q(\U6/DATA1_15 ), .QN(n1237) );
  DFFR_X2 \pipe5_divisor_n_reg[14]  ( .D(\U9/Z_14 ), .CK(clock), .RN(n1154), 
        .Q(\U6/DATA1_14 ), .QN(n1232) );
  DFFR_X2 \pipe4_divisor_n_reg[15]  ( .D(\U12/Z_15 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_15 ), .QN(n1236) );
  DFFR_X2 \pipe4_divisor_n_reg[14]  ( .D(\U12/Z_14 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_14 ), .QN(n1231) );
  DFFR_X2 \pipe3_divisor_n_reg[15]  ( .D(\U15/Z_15 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_15 ), .QN(n1235) );
  DFFR_X2 \pipe3_divisor_n_reg[14]  ( .D(\U15/Z_14 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_14 ), .QN(n1230) );
  DFFR_X2 \pipe2_divisor_n_reg[15]  ( .D(\U18/Z_15 ), .CK(clock), .RN(n1151), 
        .Q(\U15/DATA1_15 ), .QN(n1234) );
  DFFR_X2 \pipe2_divisor_n_reg[14]  ( .D(\U18/Z_14 ), .CK(clock), .RN(n1151), 
        .Q(\U15/DATA1_14 ), .QN(n1229) );
  DFFR_X2 \pipe1_divisor_n_reg[19]  ( .D(\U21/Z_19 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_19 ) );
  DFFR_X2 \pipe1_divisor_n_reg[18]  ( .D(\U21/Z_18 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_18 ) );
  DFFR_X2 \pipe1_divisor_n_reg[17]  ( .D(\U21/Z_17 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_17 ) );
  DFFR_X2 \pipe1_divisor_n_reg[16]  ( .D(\U21/Z_16 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_16 ) );
  DFFR_X2 \pipe1_divisor_n_reg[15]  ( .D(\U21/Z_15 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_15 ), .QN(n1233) );
  DFFR_X2 \pipe1_divisor_n_reg[14]  ( .D(\U21/Z_14 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_14 ), .QN(n1228) );
  DFFR_X2 \pipe1_divisor_n_reg[13]  ( .D(\U21/Z_13 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_13 ), .QN(n1223) );
  DFFR_X2 \pipe1_divisor_n_reg[12]  ( .D(\U21/Z_12 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_12 ), .QN(n1218) );
  DFFR_X2 \pipe6_divisor_n_reg[13]  ( .D(\U6/Z_13 ), .CK(clock), .RN(n1137), 
        .Q(n126) );
  DFFR_X2 \pipe6_divisor_n_reg[12]  ( .D(\U6/Z_12 ), .CK(clock), .RN(n1137), 
        .Q(n125) );
  DFFR_X2 \pipe6_divisor_n_reg[11]  ( .D(\U6/Z_11 ), .CK(clock), .RN(n1136), 
        .Q(n124) );
  DFFR_X2 \pipe6_divisor_n_reg[10]  ( .D(\U6/Z_10 ), .CK(clock), .RN(n1136), 
        .Q(n123) );
  DFFR_X2 \pipe6_divisor_n_reg[9]  ( .D(\U6/Z_9 ), .CK(clock), .RN(n1136), .Q(
        n122) );
  DFFR_X2 \pipe6_divisor_n_reg[8]  ( .D(\U6/Z_8 ), .CK(clock), .RN(n1136), .Q(
        n121) );
  DFFR_X2 \pipe6_divisor_n_reg[7]  ( .D(\U6/Z_7 ), .CK(clock), .RN(n1136), .Q(
        n120) );
  DFFR_X2 \pipe6_divisor_n_reg[6]  ( .D(\U6/Z_6 ), .CK(clock), .RN(n1136), .Q(
        n119) );
  DFFR_X2 \pipe6_divisor_n_reg[5]  ( .D(\U6/Z_5 ), .CK(clock), .RN(n1136), .Q(
        n118) );
  DFFR_X2 \pipe6_divisor_n_reg[1]  ( .D(\U6/Z_1 ), .CK(clock), .RN(n1136), .Q(
        n114) );
  DFFR_X2 \pipe5_divisor_n_reg[13]  ( .D(\U9/Z_13 ), .CK(clock), .RN(n1150), 
        .Q(\U6/DATA1_13 ), .QN(n1227) );
  DFFR_X2 \pipe5_divisor_n_reg[12]  ( .D(\U9/Z_12 ), .CK(clock), .RN(n1146), 
        .Q(\U6/DATA1_12 ), .QN(n1222) );
  DFFR_X2 \pipe5_divisor_n_reg[11]  ( .D(\U9/Z_11 ), .CK(clock), .RN(n1151), 
        .Q(\U6/DATA1_11 ), .QN(n1217) );
  DFFR_X2 \pipe5_divisor_n_reg[10]  ( .D(\U9/Z_10 ), .CK(clock), .RN(n1142), 
        .Q(\U6/DATA1_10 ), .QN(n1212) );
  DFFR_X2 \pipe5_divisor_n_reg[9]  ( .D(\U9/Z_9 ), .CK(clock), .RN(n1137), .Q(
        \U6/DATA1_9 ), .QN(n1207) );
  DFFR_X2 \pipe5_divisor_n_reg[8]  ( .D(\U9/Z_8 ), .CK(clock), .RN(n1136), .Q(
        \U6/DATA1_8 ), .QN(n1202) );
  DFFR_X2 \pipe5_divisor_n_reg[7]  ( .D(\U9/Z_7 ), .CK(clock), .RN(n1141), .Q(
        \U6/DATA1_7 ), .QN(n1197) );
  DFFR_X2 \pipe5_divisor_n_reg[6]  ( .D(\U9/Z_6 ), .CK(clock), .RN(n1145), .Q(
        \U6/DATA1_6 ), .QN(n1192) );
  DFFR_X2 \pipe5_divisor_n_reg[5]  ( .D(\U9/Z_5 ), .CK(clock), .RN(n1147), .Q(
        \U6/DATA1_5 ), .QN(n1187) );
  DFFR_X2 \pipe5_divisor_n_reg[4]  ( .D(\U9/Z_4 ), .CK(clock), .RN(n1140), .Q(
        \U6/DATA1_4 ), .QN(n1182) );
  DFFR_X2 \pipe5_divisor_n_reg[3]  ( .D(\U9/Z_3 ), .CK(clock), .RN(n1140), .Q(
        \U6/DATA1_3 ), .QN(n1177) );
  DFFR_X2 \pipe5_divisor_n_reg[2]  ( .D(\U9/Z_2 ), .CK(clock), .RN(n1140), .Q(
        \U6/DATA1_2 ), .QN(n1172) );
  DFFR_X2 \pipe5_divisor_n_reg[1]  ( .D(\U9/Z_1 ), .CK(clock), .RN(n1140), .Q(
        \U6/DATA1_1 ), .QN(n1167) );
  DFFR_X2 \pipe5_divisor_n_reg[0]  ( .D(\U9/Z_0 ), .CK(clock), .RN(n1140), .Q(
        \U6/DATA1_0 ), .QN(n1162) );
  DFFR_X2 \pipe4_divisor_n_reg[13]  ( .D(\U12/Z_13 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_13 ), .QN(n1226) );
  DFFR_X2 \pipe4_divisor_n_reg[12]  ( .D(\U12/Z_12 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_12 ), .QN(n1221) );
  DFFR_X2 \pipe4_divisor_n_reg[11]  ( .D(\U12/Z_11 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_11 ), .QN(n1216) );
  DFFR_X2 \pipe4_divisor_n_reg[10]  ( .D(\U12/Z_10 ), .CK(clock), .RN(n1147), 
        .Q(\U9/DATA1_10 ), .QN(n1211) );
  DFFR_X2 \pipe4_divisor_n_reg[9]  ( .D(\U12/Z_9 ), .CK(clock), .RN(n1133), 
        .Q(\U9/DATA1_9 ), .QN(n1206) );
  DFFR_X2 \pipe4_divisor_n_reg[8]  ( .D(\U12/Z_8 ), .CK(clock), .RN(n1135), 
        .Q(\U9/DATA1_8 ), .QN(n1201) );
  DFFR_X2 \pipe4_divisor_n_reg[7]  ( .D(\U12/Z_7 ), .CK(clock), .RN(n1152), 
        .Q(\U9/DATA1_7 ), .QN(n1196) );
  DFFR_X2 \pipe4_divisor_n_reg[6]  ( .D(\U12/Z_6 ), .CK(clock), .RN(n1149), 
        .Q(\U9/DATA1_6 ), .QN(n1191) );
  DFFR_X2 \pipe4_divisor_n_reg[5]  ( .D(\U12/Z_5 ), .CK(clock), .RN(n1137), 
        .Q(\U9/DATA1_5 ), .QN(n1186) );
  DFFR_X2 \pipe4_divisor_n_reg[4]  ( .D(\U12/Z_4 ), .CK(clock), .RN(n1143), 
        .Q(\U9/DATA1_4 ), .QN(n1181) );
  DFFR_X2 \pipe4_divisor_n_reg[3]  ( .D(\U12/Z_3 ), .CK(clock), .RN(n1138), 
        .Q(\U9/DATA1_3 ), .QN(n1176) );
  DFFR_X2 \pipe4_divisor_n_reg[2]  ( .D(\U12/Z_2 ), .CK(clock), .RN(n1153), 
        .Q(\U9/DATA1_2 ), .QN(n1171) );
  DFFR_X2 \pipe4_divisor_n_reg[1]  ( .D(\U12/Z_1 ), .CK(clock), .RN(n1148), 
        .Q(\U9/DATA1_1 ), .QN(n1166) );
  DFFR_X2 \pipe4_divisor_n_reg[0]  ( .D(\U12/Z_0 ), .CK(clock), .RN(n1144), 
        .Q(\U9/DATA1_0 ), .QN(n1161) );
  DFFR_X2 \pipe3_divisor_n_reg[13]  ( .D(\U15/Z_13 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_13 ), .QN(n1225) );
  DFFR_X2 \pipe3_divisor_n_reg[12]  ( .D(\U15/Z_12 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_12 ), .QN(n1220) );
  DFFR_X2 \pipe3_divisor_n_reg[11]  ( .D(\U15/Z_11 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_11 ), .QN(n1215) );
  DFFR_X2 \pipe3_divisor_n_reg[10]  ( .D(\U15/Z_10 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_10 ), .QN(n1210) );
  DFFR_X2 \pipe3_divisor_n_reg[9]  ( .D(\U15/Z_9 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_9 ), .QN(n1205) );
  DFFR_X2 \pipe3_divisor_n_reg[8]  ( .D(\U15/Z_8 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_8 ), .QN(n1200) );
  DFFR_X2 \pipe3_divisor_n_reg[7]  ( .D(\U15/Z_7 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_7 ), .QN(n1195) );
  DFFR_X2 \pipe3_divisor_n_reg[6]  ( .D(\U15/Z_6 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_6 ), .QN(n1190) );
  DFFR_X2 \pipe3_divisor_n_reg[5]  ( .D(\U15/Z_5 ), .CK(clock), .RN(n1145), 
        .Q(\U12/DATA1_5 ), .QN(n1185) );
  DFFR_X2 \pipe3_divisor_n_reg[4]  ( .D(\U15/Z_4 ), .CK(clock), .RN(n1145), 
        .Q(\U12/DATA1_4 ), .QN(n1180) );
  DFFR_X2 \pipe3_divisor_n_reg[3]  ( .D(\U15/Z_3 ), .CK(clock), .RN(n1145), 
        .Q(\U12/DATA1_3 ), .QN(n1175) );
  DFFR_X2 \pipe3_divisor_n_reg[2]  ( .D(\U15/Z_2 ), .CK(clock), .RN(n1145), 
        .Q(\U12/DATA1_2 ), .QN(n1170) );
  DFFR_X2 \pipe3_divisor_n_reg[1]  ( .D(\U15/Z_1 ), .CK(clock), .RN(n1145), 
        .Q(\U12/DATA1_1 ), .QN(n1165) );
  DFFR_X2 \pipe3_divisor_n_reg[0]  ( .D(\U15/Z_0 ), .CK(clock), .RN(n1145), 
        .Q(\U12/DATA1_0 ), .QN(n1160) );
  DFFR_X2 \pipe2_divisor_n_reg[13]  ( .D(\U18/Z_13 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_13 ), .QN(n1224) );
  DFFR_X2 \pipe2_divisor_n_reg[12]  ( .D(\U18/Z_12 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_12 ), .QN(n1219) );
  DFFR_X2 \pipe2_divisor_n_reg[11]  ( .D(\U18/Z_11 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_11 ), .QN(n1214) );
  DFFR_X2 \pipe2_divisor_n_reg[10]  ( .D(\U18/Z_10 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_10 ), .QN(n1209) );
  DFFR_X2 \pipe2_divisor_n_reg[9]  ( .D(\U18/Z_9 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_9 ), .QN(n1204) );
  DFFR_X2 \pipe2_divisor_n_reg[8]  ( .D(\U18/Z_8 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_8 ), .QN(n1199) );
  DFFR_X2 \pipe2_divisor_n_reg[7]  ( .D(\U18/Z_7 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_7 ), .QN(n1194) );
  DFFR_X2 \pipe2_divisor_n_reg[6]  ( .D(\U18/Z_6 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_6 ), .QN(n1189) );
  DFFR_X2 \pipe2_divisor_n_reg[5]  ( .D(\U18/Z_5 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_5 ), .QN(n1184) );
  DFFR_X2 \pipe2_divisor_n_reg[4]  ( .D(\U18/Z_4 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_4 ), .QN(n1179) );
  DFFR_X2 \pipe2_divisor_n_reg[3]  ( .D(\U18/Z_3 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_3 ), .QN(n1174) );
  DFFR_X2 \pipe2_divisor_n_reg[2]  ( .D(\U18/Z_2 ), .CK(clock), .RN(n1150), 
        .Q(\U15/DATA1_2 ), .QN(n1169) );
  DFFR_X2 \pipe2_divisor_n_reg[1]  ( .D(\U18/Z_1 ), .CK(clock), .RN(n1149), 
        .Q(\U15/DATA1_1 ), .QN(n1164) );
  DFFR_X2 \pipe2_divisor_n_reg[0]  ( .D(\U18/Z_0 ), .CK(clock), .RN(n1149), 
        .Q(\U15/DATA1_0 ), .QN(n1159) );
  DFFR_X2 \pipe1_divisor_n_reg[11]  ( .D(\U21/Z_11 ), .CK(clock), .RN(n1155), 
        .Q(\U18/DATA1_11 ), .QN(n1213) );
  DFFR_X2 \pipe1_divisor_n_reg[10]  ( .D(\U21/Z_10 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_10 ), .QN(n1208) );
  DFFR_X2 \pipe1_divisor_n_reg[9]  ( .D(\U21/Z_9 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_9 ), .QN(n1203) );
  DFFR_X2 \pipe1_divisor_n_reg[8]  ( .D(\U21/Z_8 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_8 ), .QN(n1198) );
  DFFR_X2 \pipe1_divisor_n_reg[7]  ( .D(\U21/Z_7 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_7 ), .QN(n1193) );
  DFFR_X2 \pipe1_divisor_n_reg[6]  ( .D(\U21/Z_6 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_6 ), .QN(n1188) );
  DFFR_X2 \pipe1_divisor_n_reg[5]  ( .D(\U21/Z_5 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_5 ), .QN(n1183) );
  DFFR_X2 \pipe1_divisor_n_reg[4]  ( .D(\U21/Z_4 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_4 ), .QN(n1178) );
  DFFR_X2 \pipe1_divisor_n_reg[3]  ( .D(\U21/Z_3 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_3 ), .QN(n1173) );
  DFFR_X2 \pipe1_divisor_n_reg[2]  ( .D(\U21/Z_2 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_2 ), .QN(n1168) );
  DFFR_X2 \pipe1_divisor_n_reg[1]  ( .D(\U21/Z_1 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_1 ), .QN(n1163) );
  DFFR_X2 \pipe1_divisor_n_reg[0]  ( .D(\U21/Z_0 ), .CK(clock), .RN(n1154), 
        .Q(\U18/DATA1_0 ), .QN(n1158) );
  DFFR_X2 \pipe1_result_reg[7]  ( .D(\U22/Z_7 ), .CK(clock), .RN(n1152), .Q(
        n815) );
  DFFR_X2 \pipe1_result_reg[6]  ( .D(\U22/Z_6 ), .CK(clock), .RN(n1152), .Q(
        n814) );
  DFFR_X2 \pipe1_result_reg[5]  ( .D(\U22/Z_5 ), .CK(clock), .RN(n1151), .Q(
        n813) );
  DFFR_X2 \pipe1_result_reg[4]  ( .D(\U22/Z_4 ), .CK(clock), .RN(n1151), .Q(
        n812) );
  DFFR_X2 \pipe1_result_reg[3]  ( .D(\U22/Z_3 ), .CK(clock), .RN(n1151), .Q(
        n811) );
  DFFR_X2 \pipe1_result_reg[2]  ( .D(\U22/Z_2 ), .CK(clock), .RN(n1151), .Q(
        n810) );
  DFFR_X2 \pipe1_q_reg[1]  ( .D(\U20/Z_1 ), .CK(clock), .RN(n1154), .Q(
        \U17/DATA1_2 ) );
  DFFR_X2 \pipe0_result_reg[7]  ( .D(\U25/Z_7 ), .CK(clock), .RN(n1140), .Q(
        n944) );
  DFFR_X2 \pipe0_result_reg[6]  ( .D(\U25/Z_6 ), .CK(clock), .RN(n1139), .Q(
        n943) );
  DFFR_X2 \pipe0_result_reg[5]  ( .D(\U25/Z_5 ), .CK(clock), .RN(n1134), .Q(
        n942) );
  DFFR_X2 \pipe0_result_reg[4]  ( .D(\U25/Z_4 ), .CK(clock), .RN(n1157), .Q(
        n941) );
  DFFR_X2 \pipe0_result_reg[3]  ( .D(\U25/Z_3 ), .CK(clock), .RN(n1155), .Q(
        n940) );
  DFFR_X2 \pipe0_result_reg[2]  ( .D(\U25/Z_2 ), .CK(clock), .RN(n1155), .Q(
        n939) );
  DFFR_X2 \pipe0_result_reg[1]  ( .D(\U25/Z_1 ), .CK(clock), .RN(n1155), .Q(
        n938) );
  DFFR_X2 StartOut_reg ( .D(n245), .CK(clock), .RN(n1135), .Q(StartOut) );
  DFFR_X2 StartOut5_reg ( .D(n383), .CK(clock), .RN(n1140), .Q(n245), .QN(
        n1093) );
  DFFR_X2 StartOut4_reg ( .D(n519), .CK(clock), .RN(n1154), .Q(n383), .QN(
        n1094) );
  DFFR_X2 StartOut3_reg ( .D(n653), .CK(clock), .RN(n1145), .Q(n519), .QN(
        n1095) );
  DFFR_X2 StartOut2_reg ( .D(n1098), .CK(clock), .RN(n1149), .Q(n653), .QN(
        n1092) );
  DFFR_X2 \pipe6_result_reg[7]  ( .D(\U7/Z_7 ), .CK(clock), .RN(n1133), .Q(
        n140) );
  DFFR_X2 \pipe6_result_reg[6]  ( .D(\U7/Z_6 ), .CK(clock), .RN(n1133), .Q(
        n139) );
  DFFR_X2 \pipe6_result_reg[5]  ( .D(\U7/Z_5 ), .CK(clock), .RN(n1133), .Q(
        n138) );
  DFFR_X2 \pipe6_result_reg[4]  ( .D(\U7/Z_4 ), .CK(clock), .RN(n1133), .Q(
        n137) );
  DFFR_X2 \pipe6_result_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .RN(n1133), .Q(
        n136) );
  DFFR_X2 \pipe6_result_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .RN(n1133), .Q(
        n135) );
  DFFR_X2 \pipe6_q_reg[6]  ( .D(\U5/Z_6 ), .CK(clock), .RN(n1135), .Q(
        \U4/DATA1_7 ) );
  DFFR_X2 \pipe6_q_reg[5]  ( .D(\U5/Z_5 ), .CK(clock), .RN(n1135), .Q(
        \U4/DATA1_6 ) );
  DFFR_X2 \pipe6_q_reg[4]  ( .D(\U5/Z_4 ), .CK(clock), .RN(n1135), .Q(
        \U4/DATA1_5 ) );
  DFFR_X2 \pipe6_q_reg[3]  ( .D(\U5/Z_3 ), .CK(clock), .RN(n1135), .Q(
        \U4/DATA1_4 ) );
  DFFR_X2 \pipe6_q_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .RN(n1135), .Q(
        \U4/DATA1_3 ) );
  DFFR_X2 \pipe6_q_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .RN(n1135), .Q(
        \U4/DATA1_2 ) );
  DFFR_X2 \pipe6_divisor_n_reg[19]  ( .D(\U6/Z_19 ), .CK(clock), .RN(n1137), 
        .Q(n132), .QN(n1240) );
  DFFR_X2 \pipe6_divisor_n_reg[18]  ( .D(\U6/Z_18 ), .CK(clock), .RN(n1137), 
        .Q(n131), .QN(n1239) );
  DFFR_X2 \pipe6_divisor_n_reg[17]  ( .D(\U6/Z_17 ), .CK(clock), .RN(n1137), 
        .Q(n130), .QN(n1238) );
  DFFR_X2 \pipe6_divisor_n_reg[16]  ( .D(\U6/Z_16 ), .CK(clock), .RN(n1137), 
        .Q(n129) );
  DFFR_X2 \pipe5_result_reg[7]  ( .D(\U10/Z_7 ), .CK(clock), .RN(n1138), .Q(
        n279) );
  DFFR_X2 \pipe5_result_reg[6]  ( .D(\U10/Z_6 ), .CK(clock), .RN(n1138), .Q(
        n278) );
  DFFR_X2 \pipe5_result_reg[5]  ( .D(\U10/Z_5 ), .CK(clock), .RN(n1138), .Q(
        n277) );
  DFFR_X2 \pipe5_result_reg[4]  ( .D(\U10/Z_4 ), .CK(clock), .RN(n1138), .Q(
        n276) );
  DFFR_X2 \pipe5_result_reg[3]  ( .D(\U10/Z_3 ), .CK(clock), .RN(n1137), .Q(
        n275) );
  DFFR_X2 \pipe5_result_reg[2]  ( .D(\U10/Z_2 ), .CK(clock), .RN(n1137), .Q(
        n274) );
  DFFR_X2 \pipe5_q_reg[5]  ( .D(\U8/Z_5 ), .CK(clock), .RN(n1140), .Q(
        \U5/DATA1_6 ) );
  DFFR_X2 \pipe5_q_reg[4]  ( .D(\U8/Z_4 ), .CK(clock), .RN(n1140), .Q(
        \U5/DATA1_5 ) );
  DFFR_X2 \pipe5_q_reg[3]  ( .D(\U8/Z_3 ), .CK(clock), .RN(n1140), .Q(
        \U5/DATA1_4 ) );
  DFFR_X2 \pipe5_q_reg[2]  ( .D(\U8/Z_2 ), .CK(clock), .RN(n1140), .Q(
        \U5/DATA1_3 ) );
  DFFR_X2 \pipe5_q_reg[1]  ( .D(\U8/Z_1 ), .CK(clock), .RN(n1140), .Q(
        \U5/DATA1_2 ) );
  DFFR_X2 \pipe5_divisor_n_reg[19]  ( .D(\U9/Z_19 ), .CK(clock), .RN(n1141), 
        .Q(\U6/DATA1_19 ) );
  DFFR_X2 \pipe5_divisor_n_reg[18]  ( .D(\U9/Z_18 ), .CK(clock), .RN(n1141), 
        .Q(\U6/DATA1_18 ) );
  DFFR_X2 \pipe5_divisor_n_reg[17]  ( .D(\U9/Z_17 ), .CK(clock), .RN(n1141), 
        .Q(\U6/DATA1_17 ) );
  DFFR_X2 \pipe5_divisor_n_reg[16]  ( .D(\U9/Z_16 ), .CK(clock), .RN(n1133), 
        .Q(\U6/DATA1_16 ) );
  DFFR_X2 \pipe4_result_reg[7]  ( .D(\U13/Z_7 ), .CK(clock), .RN(n1141), .Q(
        n416) );
  DFFR_X2 \pipe4_result_reg[6]  ( .D(\U13/Z_6 ), .CK(clock), .RN(n1141), .Q(
        n415) );
  DFFR_X2 \pipe4_result_reg[5]  ( .D(\U13/Z_5 ), .CK(clock), .RN(n1141), .Q(
        n414) );
  DFFR_X2 \pipe4_result_reg[4]  ( .D(\U13/Z_4 ), .CK(clock), .RN(n1141), .Q(
        n413) );
  DFFR_X2 \pipe4_result_reg[3]  ( .D(\U13/Z_3 ), .CK(clock), .RN(n1141), .Q(
        n412) );
  DFFR_X2 \pipe4_result_reg[2]  ( .D(\U13/Z_2 ), .CK(clock), .RN(n1141), .Q(
        n411) );
  DFFR_X2 \pipe4_q_reg[4]  ( .D(\U11/Z_4 ), .CK(clock), .RN(n1141), .Q(
        \U8/DATA1_5 ) );
  DFFR_X2 \pipe4_q_reg[3]  ( .D(\U11/Z_3 ), .CK(clock), .RN(n1150), .Q(
        \U8/DATA1_4 ) );
  DFFR_X2 \pipe4_q_reg[2]  ( .D(\U11/Z_2 ), .CK(clock), .RN(n1146), .Q(
        \U8/DATA1_3 ) );
  DFFR_X2 \pipe4_q_reg[1]  ( .D(\U11/Z_1 ), .CK(clock), .RN(n1151), .Q(
        \U8/DATA1_2 ) );
  DFFR_X2 \pipe4_divisor_n_reg[19]  ( .D(\U12/Z_19 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_19 ) );
  DFFR_X2 \pipe4_divisor_n_reg[18]  ( .D(\U12/Z_18 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_18 ) );
  DFFR_X2 \pipe4_divisor_n_reg[17]  ( .D(\U12/Z_17 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_17 ) );
  DFFR_X2 \pipe4_divisor_n_reg[16]  ( .D(\U12/Z_16 ), .CK(clock), .RN(n1142), 
        .Q(\U9/DATA1_16 ) );
  DFFR_X2 \pipe3_result_reg[7]  ( .D(\U16/Z_7 ), .CK(clock), .RN(n1143), .Q(
        n551) );
  DFFR_X2 \pipe3_result_reg[6]  ( .D(\U16/Z_6 ), .CK(clock), .RN(n1143), .Q(
        n550) );
  DFFR_X2 \pipe3_result_reg[5]  ( .D(\U16/Z_5 ), .CK(clock), .RN(n1143), .Q(
        n549) );
  DFFR_X2 \pipe3_result_reg[4]  ( .D(\U16/Z_4 ), .CK(clock), .RN(n1143), .Q(
        n548) );
  DFFR_X2 \pipe3_result_reg[3]  ( .D(\U16/Z_3 ), .CK(clock), .RN(n1143), .Q(
        n547) );
  DFFR_X2 \pipe3_result_reg[2]  ( .D(\U16/Z_2 ), .CK(clock), .RN(n1142), .Q(
        n546) );
  DFFR_X2 \pipe3_q_reg[3]  ( .D(\U14/Z_3 ), .CK(clock), .RN(n1145), .Q(
        \U11/DATA1_4 ) );
  DFFR_X2 \pipe3_q_reg[2]  ( .D(\U14/Z_2 ), .CK(clock), .RN(n1145), .Q(
        \U11/DATA1_3 ) );
  DFFR_X2 \pipe3_q_reg[1]  ( .D(\U14/Z_1 ), .CK(clock), .RN(n1145), .Q(
        \U11/DATA1_2 ) );
  DFFR_X2 \pipe3_divisor_n_reg[19]  ( .D(\U15/Z_19 ), .CK(clock), .RN(n1147), 
        .Q(\U12/DATA1_19 ) );
  DFFR_X2 \pipe3_divisor_n_reg[18]  ( .D(\U15/Z_18 ), .CK(clock), .RN(n1147), 
        .Q(\U12/DATA1_18 ) );
  DFFR_X2 \pipe3_divisor_n_reg[17]  ( .D(\U15/Z_17 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_17 ) );
  DFFR_X2 \pipe3_divisor_n_reg[16]  ( .D(\U15/Z_16 ), .CK(clock), .RN(n1146), 
        .Q(\U12/DATA1_16 ) );
  DFFR_X2 \pipe2_result_reg[7]  ( .D(\U19/Z_7 ), .CK(clock), .RN(n1147), .Q(
        n684) );
  DFFR_X2 \pipe2_result_reg[6]  ( .D(\U19/Z_6 ), .CK(clock), .RN(n1147), .Q(
        n683) );
  DFFR_X2 \pipe2_result_reg[5]  ( .D(\U19/Z_5 ), .CK(clock), .RN(n1147), .Q(
        n682) );
  DFFR_X2 \pipe2_result_reg[4]  ( .D(\U19/Z_4 ), .CK(clock), .RN(n1147), .Q(
        n681) );
  DFFR_X2 \pipe2_result_reg[3]  ( .D(\U19/Z_3 ), .CK(clock), .RN(n1147), .Q(
        n680) );
  DFFR_X2 \pipe2_result_reg[2]  ( .D(\U19/Z_2 ), .CK(clock), .RN(n1147), .Q(
        n679) );
  DFFR_X2 \pipe2_q_reg[2]  ( .D(\U17/Z_2 ), .CK(clock), .RN(n1149), .Q(
        \U14/DATA1_3 ) );
  DFFR_X2 \pipe2_q_reg[1]  ( .D(\U17/Z_1 ), .CK(clock), .RN(n1149), .Q(
        \U14/DATA1_2 ) );
  DFFR_X2 \pipe2_divisor_n_reg[19]  ( .D(\U18/Z_19 ), .CK(clock), .RN(n1151), 
        .Q(\U15/DATA1_19 ) );
  DFFR_X2 \pipe2_divisor_n_reg[18]  ( .D(\U18/Z_18 ), .CK(clock), .RN(n1151), 
        .Q(\U15/DATA1_18 ) );
  DFFR_X2 \pipe2_divisor_n_reg[17]  ( .D(\U18/Z_17 ), .CK(clock), .RN(n1151), 
        .Q(\U15/DATA1_17 ) );
  DFFR_X2 \pipe2_divisor_n_reg[16]  ( .D(\U18/Z_16 ), .CK(clock), .RN(n1151), 
        .Q(\U15/DATA1_16 ) );
  DFFR_X2 \pipe1_q_reg[0]  ( .D(\U20/Z_0 ), .CK(clock), .RN(n1153), .Q(
        \U17/DATA1_1 ) );
  DFFR_X2 \pipe6_q_reg[0]  ( .D(\U5/Z_0 ), .CK(clock), .RN(n1135), .Q(
        \U4/DATA1_1 ) );
  DFFR_X2 \pipe5_q_reg[0]  ( .D(\U8/Z_0 ), .CK(clock), .RN(n1140), .Q(
        \U5/DATA1_1 ) );
  DFFR_X2 \pipe4_q_reg[0]  ( .D(\U11/Z_0 ), .CK(clock), .RN(n1142), .Q(
        \U8/DATA1_1 ) );
  DFFR_X2 \pipe3_q_reg[0]  ( .D(\U14/Z_0 ), .CK(clock), .RN(n1145), .Q(
        \U11/DATA1_1 ) );
  DFFR_X2 \pipe2_q_reg[0]  ( .D(\U17/Z_0 ), .CK(clock), .RN(n1149), .Q(
        \U14/DATA1_1 ) );
  DFFR_X2 \pipe1_result_reg[14]  ( .D(\U22/Z_14 ), .CK(clock), .RN(n1152), .Q(
        n822) );
  DFFR_X2 \pipe1_result_reg[13]  ( .D(\U22/Z_13 ), .CK(clock), .RN(n1152), .Q(
        n821) );
  DFFR_X2 \pipe1_result_reg[10]  ( .D(\U22/Z_10 ), .CK(clock), .RN(n1152), .Q(
        n818) );
  DFFR_X2 \pipe1_result_reg[9]  ( .D(\U22/Z_9 ), .CK(clock), .RN(n1152), .Q(
        n817) );
  DFFR_X2 \pipe1_result_reg[18]  ( .D(\U22/Z_18 ), .CK(clock), .RN(n1153), .Q(
        n826) );
  DFFR_X2 \pipe1_result_reg[15]  ( .D(\U22/Z_15 ), .CK(clock), .RN(n1152), .Q(
        n823) );
  DFFR_X2 \pipe6_divisor_n_reg[4]  ( .D(\U6/Z_4 ), .CK(clock), .RN(n1136), .Q(
        n117) );
  DFFR_X2 \pipe6_divisor_n_reg[3]  ( .D(\U6/Z_3 ), .CK(clock), .RN(n1136), .Q(
        n116) );
  DFFR_X2 \pipe6_divisor_n_reg[2]  ( .D(\U6/Z_2 ), .CK(clock), .RN(n1136), .Q(
        n115) );
  DFFR_X2 \pipe0_q_reg[0]  ( .D(\U23/Z_0 ), .CK(clock), .RN(n1157), .Q(
        \U20/DATA1_1 ) );
  DFFR_X2 \pipe0_result_reg[12]  ( .D(\U25/Z_12 ), .CK(clock), .RN(n1156), .Q(
        n949) );
  DFFR_X2 \pipe0_result_reg[17]  ( .D(\U25/Z_17 ), .CK(clock), .RN(reset_n), 
        .Q(n954) );
  DFFR_X2 \pipe0_result_reg[13]  ( .D(\U25/Z_13 ), .CK(clock), .RN(n1151), .Q(
        n950) );
  DFFR_X2 \pipe0_result_reg[11]  ( .D(\U25/Z_11 ), .CK(clock), .RN(n1142), .Q(
        n948) );
  DFFR_X2 \pipe6_result_reg[8]  ( .D(\U7/Z_8 ), .CK(clock), .RN(n1133), .Q(
        n141) );
  DFFR_X2 \pipe6_result_reg[11]  ( .D(\U7/Z_11 ), .CK(clock), .RN(n1133), .Q(
        n144) );
  DFFR_X2 \pipe0_result_reg[10]  ( .D(\U25/Z_10 ), .CK(clock), .RN(n1137), .Q(
        n947) );
  DFFR_X2 \pipe0_result_reg[9]  ( .D(\U25/Z_9 ), .CK(clock), .RN(n1141), .Q(
        n946) );
  DFFR_X2 \pipe0_result_reg[8]  ( .D(\U25/Z_8 ), .CK(clock), .RN(n1147), .Q(
        n945) );
  DFFR_X2 \pipe0_result_reg[18]  ( .D(\U25/Z_18 ), .CK(clock), .RN(n1156), .Q(
        n955) );
  DFFR_X2 \pipe0_result_reg[16]  ( .D(\U25/Z_16 ), .CK(clock), .RN(n1156), .Q(
        n953) );
  DFFR_X2 \pipe0_result_reg[15]  ( .D(\U25/Z_15 ), .CK(clock), .RN(n1156), .Q(
        n952) );
  DFFR_X2 \pipe0_result_reg[14]  ( .D(\U25/Z_14 ), .CK(clock), .RN(n1133), .Q(
        n951) );
  DFFR_X2 \pipe0_result_reg[19]  ( .D(\U25/Z_19 ), .CK(clock), .RN(n1156), .Q(
        n956) );
  DFFR_X2 \pipe0_result_reg[27]  ( .D(\U25/Z_27 ), .CK(clock), .RN(n1157), .Q(
        n964) );
  DFFR_X2 \pipe0_result_reg[26]  ( .D(\U25/Z_26 ), .CK(clock), .RN(n1156), .Q(
        n963) );
  DFFR_X2 \pipe0_result_reg[25]  ( .D(\U25/Z_25 ), .CK(clock), .RN(n1156), .Q(
        n962) );
  DFFR_X2 \pipe0_result_reg[24]  ( .D(\U25/Z_24 ), .CK(clock), .RN(n1156), .Q(
        n961) );
  DFFR_X2 \pipe0_result_reg[23]  ( .D(\U25/Z_23 ), .CK(clock), .RN(n1156), .Q(
        n960) );
  DFFR_X2 \pipe0_result_reg[22]  ( .D(\U25/Z_22 ), .CK(clock), .RN(n1156), .Q(
        n959) );
  INV_X4 U23 ( .A(divisor[6]), .ZN(n1257) );
  AND2_X4 U24 ( .A1(\U4/DATA1_0 ), .A2(n41), .ZN(\U4/Z_0 ) );
  INV_X4 U25 ( .A(divisor[10]), .ZN(n1253) );
  INV_X1 U26 ( .A(n1254), .ZN(n1119) );
  INV_X4 U27 ( .A(n1119), .ZN(n1120) );
  INV_X4 U28 ( .A(divisor[15]), .ZN(n1248) );
  INV_X4 U29 ( .A(divisor[19]), .ZN(n1121) );
  INV_X1 U30 ( .A(n1250), .ZN(n1122) );
  INV_X4 U31 ( .A(n1122), .ZN(n1123) );
  INV_X1 U32 ( .A(n1259), .ZN(n1124) );
  INV_X4 U33 ( .A(n1124), .ZN(n1125) );
  INV_X4 U34 ( .A(divisor[17]), .ZN(n1126) );
  INV_X4 U35 ( .A(divisor[9]), .ZN(n1254) );
  INV_X4 U36 ( .A(divisor[1]), .ZN(n1262) );
  INV_X4 U37 ( .A(divisor[18]), .ZN(n1127) );
  OR3_X1 U38 ( .A1(n115), .A2(n116), .A3(n117), .ZN(n1128) );
  OR3_X4 U39 ( .A1(n114), .A2(n113), .A3(n1128), .ZN(n1244) );
  OR3_X4 U40 ( .A1(n124), .A2(n123), .A3(n1129), .ZN(n1242) );
  BUF_X4 U41 ( .A(reset_n), .Z(n1136) );
  BUF_X4 U42 ( .A(reset_n), .Z(n1134) );
  BUF_X4 U43 ( .A(reset_n), .Z(n1135) );
  BUF_X4 U44 ( .A(reset_n), .Z(n1138) );
  BUF_X4 U45 ( .A(reset_n), .Z(n1139) );
  BUF_X4 U46 ( .A(reset_n), .Z(n1140) );
  BUF_X4 U47 ( .A(reset_n), .Z(n1143) );
  BUF_X4 U48 ( .A(reset_n), .Z(n1144) );
  BUF_X4 U49 ( .A(reset_n), .Z(n1145) );
  BUF_X4 U50 ( .A(reset_n), .Z(n1146) );
  BUF_X4 U51 ( .A(reset_n), .Z(n1148) );
  BUF_X4 U52 ( .A(reset_n), .Z(n1149) );
  BUF_X4 U53 ( .A(reset_n), .Z(n1150) );
  BUF_X4 U54 ( .A(reset_n), .Z(n1152) );
  BUF_X4 U55 ( .A(reset_n), .Z(n1153) );
  BUF_X4 U60 ( .A(reset_n), .Z(n1154) );
  BUF_X4 U61 ( .A(reset_n), .Z(n1157) );
  BUF_X4 U62 ( .A(reset_n), .Z(n1156) );
  BUF_X4 U63 ( .A(reset_n), .Z(n1133) );
  BUF_X4 U64 ( .A(reset_n), .Z(n1137) );
  BUF_X4 U65 ( .A(reset_n), .Z(n1141) );
  BUF_X4 U66 ( .A(reset_n), .Z(n1142) );
  BUF_X4 U67 ( .A(reset_n), .Z(n1147) );
  BUF_X4 U72 ( .A(reset_n), .Z(n1151) );
  BUF_X4 U73 ( .A(reset_n), .Z(n1155) );
  INV_X4 U74 ( .A(n1132), .ZN(n1131) );
  OR3_X4 U75 ( .A1(n125), .A2(n126), .A3(n127), .ZN(n1129) );
  OR3_X1 U76 ( .A1(n122), .A2(n121), .A3(n120), .ZN(n1243) );
  INV_X4 U81 ( .A(start), .ZN(n1132) );
  AND2_X4 U90 ( .A1(\U23/DATA1_0 ), .A2(n1131), .ZN(\U23/Z_0 ) );
  INV_X4 U91 ( .A(divisor[0]), .ZN(n1263) );
  NOR2_X2 U92 ( .A1(n1130), .A2(n1099), .ZN(\U21/Z_0 ) );
  NOR2_X2 U93 ( .A1(n1096), .A2(n1158), .ZN(\U18/Z_0 ) );
  NOR2_X2 U94 ( .A1(n1092), .A2(n1159), .ZN(\U15/Z_0 ) );
  NOR2_X2 U95 ( .A1(n1095), .A2(n1160), .ZN(\U12/Z_0 ) );
  NOR2_X2 U96 ( .A1(n1094), .A2(n1161), .ZN(\U9/Z_0 ) );
  NOR2_X2 U97 ( .A1(n1093), .A2(n1162), .ZN(\U6/Z_0 ) );
  NOR2_X2 U98 ( .A1(n1130), .A2(n1100), .ZN(\U21/Z_1 ) );
  NOR2_X2 U99 ( .A1(n1096), .A2(n1163), .ZN(\U18/Z_1 ) );
  NOR2_X2 U101 ( .A1(n1092), .A2(n1164), .ZN(\U15/Z_1 ) );
  NOR2_X2 U102 ( .A1(n1095), .A2(n1165), .ZN(\U12/Z_1 ) );
  NOR2_X2 U103 ( .A1(n1094), .A2(n1166), .ZN(\U9/Z_1 ) );
  NOR2_X2 U104 ( .A1(n1093), .A2(n1167), .ZN(\U6/Z_1 ) );
  INV_X4 U105 ( .A(divisor[2]), .ZN(n1261) );
  NOR2_X2 U106 ( .A1(n1130), .A2(n1101), .ZN(\U21/Z_2 ) );
  NOR2_X2 U107 ( .A1(n1096), .A2(n1168), .ZN(\U18/Z_2 ) );
  NOR2_X2 U108 ( .A1(n1092), .A2(n1169), .ZN(\U15/Z_2 ) );
  NOR2_X2 U109 ( .A1(n1095), .A2(n1170), .ZN(\U12/Z_2 ) );
  NOR2_X2 U114 ( .A1(n1094), .A2(n1171), .ZN(\U9/Z_2 ) );
  NOR2_X2 U115 ( .A1(n1093), .A2(n1172), .ZN(\U6/Z_2 ) );
  INV_X4 U116 ( .A(divisor[3]), .ZN(n1260) );
  NOR2_X2 U117 ( .A1(n1130), .A2(n1102), .ZN(\U21/Z_3 ) );
  NOR2_X2 U118 ( .A1(n1096), .A2(n1173), .ZN(\U18/Z_3 ) );
  NOR2_X2 U119 ( .A1(n1092), .A2(n1174), .ZN(\U15/Z_3 ) );
  NOR2_X2 U120 ( .A1(n1095), .A2(n1175), .ZN(\U12/Z_3 ) );
  NOR2_X2 U121 ( .A1(n1094), .A2(n1176), .ZN(\U9/Z_3 ) );
  NOR2_X2 U127 ( .A1(n1093), .A2(n1177), .ZN(\U6/Z_3 ) );
  INV_X4 U128 ( .A(divisor[4]), .ZN(n1259) );
  NOR2_X2 U135 ( .A1(n1130), .A2(n1103), .ZN(\U21/Z_4 ) );
  NOR2_X2 U136 ( .A1(n1096), .A2(n1178), .ZN(\U18/Z_4 ) );
  NOR2_X2 U137 ( .A1(n1092), .A2(n1179), .ZN(\U15/Z_4 ) );
  NOR2_X2 U138 ( .A1(n1095), .A2(n1180), .ZN(\U12/Z_4 ) );
  NOR2_X2 U139 ( .A1(n1094), .A2(n1181), .ZN(\U9/Z_4 ) );
  NOR2_X2 U140 ( .A1(n1093), .A2(n1182), .ZN(\U6/Z_4 ) );
  INV_X4 U141 ( .A(divisor[5]), .ZN(n1258) );
  NOR2_X2 U142 ( .A1(n1130), .A2(n1104), .ZN(\U21/Z_5 ) );
  NOR2_X2 U143 ( .A1(n1096), .A2(n1183), .ZN(\U18/Z_5 ) );
  NOR2_X2 U148 ( .A1(n1092), .A2(n1184), .ZN(\U15/Z_5 ) );
  NOR2_X2 U149 ( .A1(n1095), .A2(n1185), .ZN(\U12/Z_5 ) );
  NOR2_X2 U150 ( .A1(n1094), .A2(n1186), .ZN(\U9/Z_5 ) );
  NOR2_X2 U151 ( .A1(n1093), .A2(n1187), .ZN(\U6/Z_5 ) );
  NOR2_X2 U152 ( .A1(n1130), .A2(n1105), .ZN(\U21/Z_6 ) );
  NOR2_X2 U153 ( .A1(n1096), .A2(n1188), .ZN(\U18/Z_6 ) );
  NOR2_X2 U154 ( .A1(n1092), .A2(n1189), .ZN(\U15/Z_6 ) );
  NOR2_X2 U155 ( .A1(n1095), .A2(n1190), .ZN(\U12/Z_6 ) );
  NOR2_X2 U157 ( .A1(n1094), .A2(n1191), .ZN(\U9/Z_6 ) );
  NOR2_X2 U158 ( .A1(n1093), .A2(n1192), .ZN(\U6/Z_6 ) );
  INV_X4 U159 ( .A(divisor[7]), .ZN(n1256) );
  NOR2_X2 U160 ( .A1(n1130), .A2(n1106), .ZN(\U21/Z_7 ) );
  NOR2_X2 U161 ( .A1(n1096), .A2(n1193), .ZN(\U18/Z_7 ) );
  NOR2_X2 U162 ( .A1(n1092), .A2(n1194), .ZN(\U15/Z_7 ) );
  NOR2_X2 U163 ( .A1(n1095), .A2(n1195), .ZN(\U12/Z_7 ) );
  NOR2_X2 U164 ( .A1(n1094), .A2(n1196), .ZN(\U9/Z_7 ) );
  NOR2_X2 U165 ( .A1(n1093), .A2(n1197), .ZN(\U6/Z_7 ) );
  INV_X4 U166 ( .A(divisor[8]), .ZN(n1255) );
  NOR2_X2 U168 ( .A1(n1130), .A2(n1107), .ZN(\U21/Z_8 ) );
  NOR2_X2 U169 ( .A1(n1096), .A2(n1198), .ZN(\U18/Z_8 ) );
  NOR2_X2 U170 ( .A1(n1092), .A2(n1199), .ZN(\U15/Z_8 ) );
  NOR2_X2 U171 ( .A1(n1095), .A2(n1200), .ZN(\U12/Z_8 ) );
  NOR2_X2 U172 ( .A1(n1094), .A2(n1201), .ZN(\U9/Z_8 ) );
  NOR2_X2 U177 ( .A1(n1093), .A2(n1202), .ZN(\U6/Z_8 ) );
  NOR2_X2 U178 ( .A1(n1130), .A2(n1108), .ZN(\U21/Z_9 ) );
  NOR2_X2 U179 ( .A1(n1096), .A2(n1203), .ZN(\U18/Z_9 ) );
  NOR2_X2 U180 ( .A1(n1092), .A2(n1204), .ZN(\U15/Z_9 ) );
  NOR2_X2 U181 ( .A1(n1095), .A2(n1205), .ZN(\U12/Z_9 ) );
  NOR2_X2 U182 ( .A1(n1094), .A2(n1206), .ZN(\U9/Z_9 ) );
  NOR2_X2 U183 ( .A1(n1093), .A2(n1207), .ZN(\U6/Z_9 ) );
  NOR2_X2 U184 ( .A1(n1130), .A2(n1109), .ZN(\U21/Z_10 ) );
  NOR2_X2 U186 ( .A1(n1096), .A2(n1208), .ZN(\U18/Z_10 ) );
  NOR2_X2 U187 ( .A1(n1092), .A2(n1209), .ZN(\U15/Z_10 ) );
  NOR2_X2 U188 ( .A1(n1095), .A2(n1210), .ZN(\U12/Z_10 ) );
  NOR2_X2 U189 ( .A1(n1094), .A2(n1211), .ZN(\U9/Z_10 ) );
  NOR2_X2 U190 ( .A1(n1093), .A2(n1212), .ZN(\U6/Z_10 ) );
  INV_X4 U191 ( .A(divisor[11]), .ZN(n1252) );
  NOR2_X2 U192 ( .A1(n1130), .A2(n1110), .ZN(\U21/Z_11 ) );
  NOR2_X2 U193 ( .A1(n1096), .A2(n1213), .ZN(\U18/Z_11 ) );
  NOR2_X2 U194 ( .A1(n1092), .A2(n1214), .ZN(\U15/Z_11 ) );
  NOR2_X2 U195 ( .A1(n1095), .A2(n1215), .ZN(\U12/Z_11 ) );
  NOR2_X2 U197 ( .A1(n1094), .A2(n1216), .ZN(\U9/Z_11 ) );
  NOR2_X2 U198 ( .A1(n1093), .A2(n1217), .ZN(\U6/Z_11 ) );
  INV_X4 U199 ( .A(divisor[12]), .ZN(n1251) );
  NOR2_X2 U200 ( .A1(n1130), .A2(n1111), .ZN(\U21/Z_12 ) );
  NOR2_X2 U201 ( .A1(n1096), .A2(n1218), .ZN(\U18/Z_12 ) );
  NOR2_X2 U202 ( .A1(n1092), .A2(n1219), .ZN(\U15/Z_12 ) );
  NOR2_X2 U203 ( .A1(n1095), .A2(n1220), .ZN(\U12/Z_12 ) );
  NOR2_X2 U204 ( .A1(n1094), .A2(n1221), .ZN(\U9/Z_12 ) );
  NOR2_X2 U205 ( .A1(n1093), .A2(n1222), .ZN(\U6/Z_12 ) );
  INV_X4 U206 ( .A(divisor[13]), .ZN(n1250) );
  NOR2_X2 U207 ( .A1(n1130), .A2(n1112), .ZN(\U21/Z_13 ) );
  NOR2_X2 U208 ( .A1(n1096), .A2(n1223), .ZN(\U18/Z_13 ) );
  NOR2_X2 U209 ( .A1(n1092), .A2(n1224), .ZN(\U15/Z_13 ) );
  NOR2_X2 U210 ( .A1(n1095), .A2(n1225), .ZN(\U12/Z_13 ) );
  NOR2_X2 U211 ( .A1(n1094), .A2(n1226), .ZN(\U9/Z_13 ) );
  NOR2_X2 U212 ( .A1(n1093), .A2(n1227), .ZN(\U6/Z_13 ) );
  INV_X4 U213 ( .A(divisor[14]), .ZN(n1249) );
  NOR2_X2 U214 ( .A1(n1130), .A2(n1113), .ZN(\U21/Z_14 ) );
  NOR2_X2 U215 ( .A1(n1096), .A2(n1228), .ZN(\U18/Z_14 ) );
  NOR2_X2 U216 ( .A1(n1092), .A2(n1229), .ZN(\U15/Z_14 ) );
  NOR2_X2 U217 ( .A1(n1095), .A2(n1230), .ZN(\U12/Z_14 ) );
  NOR2_X2 U218 ( .A1(n1094), .A2(n1231), .ZN(\U9/Z_14 ) );
  NOR2_X2 U219 ( .A1(n1093), .A2(n1232), .ZN(\U6/Z_14 ) );
  NOR2_X2 U220 ( .A1(n1130), .A2(n1114), .ZN(\U21/Z_15 ) );
  NOR2_X2 U221 ( .A1(n1096), .A2(n1233), .ZN(\U18/Z_15 ) );
  NOR2_X2 U222 ( .A1(n1092), .A2(n1234), .ZN(\U15/Z_15 ) );
  NOR2_X2 U227 ( .A1(n1095), .A2(n1235), .ZN(\U12/Z_15 ) );
  NOR2_X2 U228 ( .A1(n1094), .A2(n1236), .ZN(\U9/Z_15 ) );
  NOR2_X2 U229 ( .A1(n1093), .A2(n1237), .ZN(\U6/Z_15 ) );
  AND2_X1 U230 ( .A1(\U7/DATA1_7 ), .A2(n245), .ZN(\U7/Z_7 ) );
  AND2_X1 U231 ( .A1(\U7/DATA1_8 ), .A2(n245), .ZN(\U7/Z_8 ) );
  AND2_X1 U232 ( .A1(\U7/DATA1_9 ), .A2(n245), .ZN(\U7/Z_9 ) );
  AND2_X1 U233 ( .A1(\U7/DATA1_10 ), .A2(n245), .ZN(\U7/Z_10 ) );
  AND2_X1 U234 ( .A1(\U7/DATA1_11 ), .A2(n245), .ZN(\U7/Z_11 ) );
  AND2_X1 U236 ( .A1(\U7/DATA1_12 ), .A2(n245), .ZN(\U7/Z_12 ) );
  AND2_X1 U237 ( .A1(\U7/DATA1_13 ), .A2(n245), .ZN(\U7/Z_13 ) );
  AND2_X1 U238 ( .A1(\U7/DATA1_14 ), .A2(n245), .ZN(\U7/Z_14 ) );
  AND2_X1 U239 ( .A1(\U7/DATA1_15 ), .A2(n245), .ZN(\U7/Z_15 ) );
  AND2_X1 U240 ( .A1(\U7/DATA1_16 ), .A2(n245), .ZN(\U7/Z_16 ) );
  AND2_X1 U241 ( .A1(\U7/DATA1_17 ), .A2(n245), .ZN(\U7/Z_17 ) );
  AND2_X1 U242 ( .A1(\U7/DATA1_18 ), .A2(n245), .ZN(\U7/Z_18 ) );
  AND2_X1 U243 ( .A1(\U7/DATA1_19 ), .A2(n245), .ZN(\U7/Z_19 ) );
  AND2_X1 U244 ( .A1(\U7/DATA1_20 ), .A2(n245), .ZN(\U7/Z_20 ) );
  AND2_X1 U245 ( .A1(\U7/DATA1_21 ), .A2(n245), .ZN(\U7/Z_21 ) );
  AND2_X1 U247 ( .A1(\U7/DATA1_22 ), .A2(n245), .ZN(\U7/Z_22 ) );
  AND2_X1 U248 ( .A1(\U7/DATA1_23 ), .A2(n245), .ZN(\U7/Z_23 ) );
  AND2_X1 U249 ( .A1(\U7/DATA1_24 ), .A2(n245), .ZN(\U7/Z_24 ) );
  AND2_X1 U250 ( .A1(\U7/DATA1_25 ), .A2(n245), .ZN(\U7/Z_25 ) );
  AND2_X1 U251 ( .A1(\U7/DATA1_26 ), .A2(n245), .ZN(\U7/Z_26 ) );
  AND2_X1 U252 ( .A1(\U7/DATA1_27 ), .A2(n245), .ZN(\U7/Z_27 ) );
  AND2_X1 U253 ( .A1(\U10/DATA1_7 ), .A2(n383), .ZN(\U10/Z_7 ) );
  AND2_X1 U254 ( .A1(\U10/DATA1_8 ), .A2(n383), .ZN(\U10/Z_8 ) );
  AND2_X1 U255 ( .A1(\U10/DATA1_9 ), .A2(n383), .ZN(\U10/Z_9 ) );
  AND2_X1 U260 ( .A1(\U10/DATA1_10 ), .A2(n383), .ZN(\U10/Z_10 ) );
  AND2_X1 U261 ( .A1(\U10/DATA1_11 ), .A2(n383), .ZN(\U10/Z_11 ) );
  AND2_X1 U262 ( .A1(\U10/DATA1_12 ), .A2(n383), .ZN(\U10/Z_12 ) );
  AND2_X1 U263 ( .A1(\U10/DATA1_13 ), .A2(n383), .ZN(\U10/Z_13 ) );
  AND2_X1 U264 ( .A1(\U10/DATA1_14 ), .A2(n383), .ZN(\U10/Z_14 ) );
  AND2_X1 U265 ( .A1(\U10/DATA1_15 ), .A2(n383), .ZN(\U10/Z_15 ) );
  AND2_X1 U266 ( .A1(\U10/DATA1_16 ), .A2(n383), .ZN(\U10/Z_16 ) );
  AND2_X1 U267 ( .A1(\U10/DATA1_17 ), .A2(n383), .ZN(\U10/Z_17 ) );
  AND2_X1 U269 ( .A1(\U10/DATA1_18 ), .A2(n383), .ZN(\U10/Z_18 ) );
  AND2_X1 U270 ( .A1(\U10/DATA1_19 ), .A2(n383), .ZN(\U10/Z_19 ) );
  AND2_X1 U271 ( .A1(\U10/DATA1_20 ), .A2(n383), .ZN(\U10/Z_20 ) );
  AND2_X1 U272 ( .A1(\U10/DATA1_21 ), .A2(n383), .ZN(\U10/Z_21 ) );
  AND2_X1 U273 ( .A1(\U10/DATA1_22 ), .A2(n383), .ZN(\U10/Z_22 ) );
  AND2_X1 U278 ( .A1(\U10/DATA1_23 ), .A2(n383), .ZN(\U10/Z_23 ) );
  AND2_X1 U279 ( .A1(\U10/DATA1_24 ), .A2(n383), .ZN(\U10/Z_24 ) );
  AND2_X1 U280 ( .A1(\U10/DATA1_25 ), .A2(n383), .ZN(\U10/Z_25 ) );
  AND2_X1 U281 ( .A1(\U10/DATA1_26 ), .A2(n383), .ZN(\U10/Z_26 ) );
  AND2_X1 U282 ( .A1(\U10/DATA1_27 ), .A2(n383), .ZN(\U10/Z_27 ) );
  AND2_X1 U283 ( .A1(\U13/DATA1_7 ), .A2(n519), .ZN(\U13/Z_7 ) );
  AND2_X1 U284 ( .A1(\U13/DATA1_8 ), .A2(n519), .ZN(\U13/Z_8 ) );
  AND2_X1 U285 ( .A1(\U13/DATA1_9 ), .A2(n519), .ZN(\U13/Z_9 ) );
  AND2_X1 U287 ( .A1(\U13/DATA1_10 ), .A2(n519), .ZN(\U13/Z_10 ) );
  AND2_X1 U288 ( .A1(\U13/DATA1_11 ), .A2(n519), .ZN(\U13/Z_11 ) );
  AND2_X1 U289 ( .A1(\U13/DATA1_12 ), .A2(n519), .ZN(\U13/Z_12 ) );
  AND2_X1 U290 ( .A1(\U13/DATA1_13 ), .A2(n519), .ZN(\U13/Z_13 ) );
  AND2_X1 U291 ( .A1(\U13/DATA1_14 ), .A2(n519), .ZN(\U13/Z_14 ) );
  AND2_X1 U292 ( .A1(\U13/DATA1_15 ), .A2(n519), .ZN(\U13/Z_15 ) );
  AND2_X1 U293 ( .A1(\U13/DATA1_16 ), .A2(n519), .ZN(\U13/Z_16 ) );
  AND2_X1 U294 ( .A1(\U13/DATA1_17 ), .A2(n519), .ZN(\U13/Z_17 ) );
  AND2_X1 U295 ( .A1(\U13/DATA1_18 ), .A2(n519), .ZN(\U13/Z_18 ) );
  AND2_X1 U296 ( .A1(\U13/DATA1_19 ), .A2(n519), .ZN(\U13/Z_19 ) );
  AND2_X1 U298 ( .A1(\U13/DATA1_20 ), .A2(n519), .ZN(\U13/Z_20 ) );
  AND2_X1 U299 ( .A1(\U13/DATA1_21 ), .A2(n519), .ZN(\U13/Z_21 ) );
  AND2_X1 U300 ( .A1(\U13/DATA1_22 ), .A2(n519), .ZN(\U13/Z_22 ) );
  AND2_X1 U301 ( .A1(\U13/DATA1_23 ), .A2(n519), .ZN(\U13/Z_23 ) );
  AND2_X1 U302 ( .A1(\U13/DATA1_24 ), .A2(n519), .ZN(\U13/Z_24 ) );
  AND2_X1 U303 ( .A1(\U13/DATA1_25 ), .A2(n519), .ZN(\U13/Z_25 ) );
  AND2_X1 U304 ( .A1(\U13/DATA1_26 ), .A2(n519), .ZN(\U13/Z_26 ) );
  AND2_X1 U305 ( .A1(\U13/DATA1_27 ), .A2(n519), .ZN(\U13/Z_27 ) );
  AND2_X1 U306 ( .A1(\U16/DATA1_7 ), .A2(n653), .ZN(\U16/Z_7 ) );
  AND2_X1 U311 ( .A1(\U16/DATA1_8 ), .A2(n653), .ZN(\U16/Z_8 ) );
  AND2_X1 U312 ( .A1(\U16/DATA1_9 ), .A2(n653), .ZN(\U16/Z_9 ) );
  AND2_X1 U313 ( .A1(\U16/DATA1_10 ), .A2(n653), .ZN(\U16/Z_10 ) );
  AND2_X1 U314 ( .A1(\U16/DATA1_11 ), .A2(n653), .ZN(\U16/Z_11 ) );
  AND2_X1 U315 ( .A1(\U16/DATA1_12 ), .A2(n653), .ZN(\U16/Z_12 ) );
  AND2_X1 U316 ( .A1(\U16/DATA1_13 ), .A2(n653), .ZN(\U16/Z_13 ) );
  AND2_X1 U317 ( .A1(\U16/DATA1_14 ), .A2(n653), .ZN(\U16/Z_14 ) );
  AND2_X1 U318 ( .A1(\U16/DATA1_15 ), .A2(n653), .ZN(\U16/Z_15 ) );
  AND2_X1 U321 ( .A1(\U16/DATA1_16 ), .A2(n653), .ZN(\U16/Z_16 ) );
  AND2_X1 U322 ( .A1(\U16/DATA1_17 ), .A2(n653), .ZN(\U16/Z_17 ) );
  AND2_X1 U323 ( .A1(\U16/DATA1_18 ), .A2(n653), .ZN(\U16/Z_18 ) );
  AND2_X1 U324 ( .A1(\U16/DATA1_19 ), .A2(n653), .ZN(\U16/Z_19 ) );
  AND2_X1 U325 ( .A1(\U16/DATA1_20 ), .A2(n653), .ZN(\U16/Z_20 ) );
  AND2_X1 U330 ( .A1(\U16/DATA1_21 ), .A2(n653), .ZN(\U16/Z_21 ) );
  AND2_X1 U331 ( .A1(\U16/DATA1_22 ), .A2(n653), .ZN(\U16/Z_22 ) );
  AND2_X1 U332 ( .A1(\U16/DATA1_23 ), .A2(n653), .ZN(\U16/Z_23 ) );
  AND2_X1 U333 ( .A1(\U16/DATA1_24 ), .A2(n653), .ZN(\U16/Z_24 ) );
  AND2_X1 U334 ( .A1(\U16/DATA1_25 ), .A2(n653), .ZN(\U16/Z_25 ) );
  AND2_X1 U335 ( .A1(\U16/DATA1_26 ), .A2(n653), .ZN(\U16/Z_26 ) );
  AND2_X1 U336 ( .A1(\U16/DATA1_27 ), .A2(n653), .ZN(\U16/Z_27 ) );
  AND2_X1 U337 ( .A1(\U19/DATA1_7 ), .A2(n1098), .ZN(\U19/Z_7 ) );
  AND2_X1 U339 ( .A1(\U19/DATA1_8 ), .A2(n1098), .ZN(\U19/Z_8 ) );
  AND2_X1 U340 ( .A1(\U19/DATA1_9 ), .A2(n1098), .ZN(\U19/Z_9 ) );
  AND2_X1 U341 ( .A1(\U19/DATA1_10 ), .A2(n1098), .ZN(\U19/Z_10 ) );
  AND2_X1 U342 ( .A1(\U19/DATA1_11 ), .A2(n1098), .ZN(\U19/Z_11 ) );
  AND2_X1 U343 ( .A1(\U19/DATA1_12 ), .A2(n1098), .ZN(\U19/Z_12 ) );
  AND2_X1 U344 ( .A1(\U19/DATA1_13 ), .A2(n1098), .ZN(\U19/Z_13 ) );
  AND2_X1 U345 ( .A1(\U19/DATA1_14 ), .A2(n1098), .ZN(\U19/Z_14 ) );
  AND2_X1 U346 ( .A1(\U19/DATA1_15 ), .A2(n1098), .ZN(\U19/Z_15 ) );
  AND2_X1 U347 ( .A1(\U19/DATA1_16 ), .A2(n1098), .ZN(\U19/Z_16 ) );
  AND2_X1 U348 ( .A1(\U19/DATA1_17 ), .A2(n1098), .ZN(\U19/Z_17 ) );
  AND2_X1 U350 ( .A1(\U19/DATA1_18 ), .A2(n1098), .ZN(\U19/Z_18 ) );
  AND2_X1 U351 ( .A1(\U19/DATA1_19 ), .A2(n1098), .ZN(\U19/Z_19 ) );
  AND2_X1 U352 ( .A1(\U19/DATA1_20 ), .A2(n1098), .ZN(\U19/Z_20 ) );
  AND2_X1 U353 ( .A1(\U19/DATA1_21 ), .A2(n1098), .ZN(\U19/Z_21 ) );
  AND2_X1 U354 ( .A1(\U19/DATA1_22 ), .A2(n1098), .ZN(\U19/Z_22 ) );
  AND2_X1 U355 ( .A1(\U19/DATA1_23 ), .A2(n1098), .ZN(\U19/Z_23 ) );
  AND2_X1 U356 ( .A1(\U19/DATA1_24 ), .A2(n1098), .ZN(\U19/Z_24 ) );
  AND2_X1 U357 ( .A1(\U19/DATA1_25 ), .A2(n1098), .ZN(\U19/Z_25 ) );
  AND2_X1 U358 ( .A1(\U19/DATA1_26 ), .A2(n1098), .ZN(\U19/Z_26 ) );
  AND2_X1 U363 ( .A1(\U19/DATA1_27 ), .A2(n1098), .ZN(\U19/Z_27 ) );
  AND2_X1 U364 ( .A1(\U22/DATA1_7 ), .A2(n915), .ZN(\U22/Z_7 ) );
  AND2_X1 U365 ( .A1(\U22/DATA1_8 ), .A2(n915), .ZN(\U22/Z_8 ) );
  AND2_X1 U366 ( .A1(\U22/DATA1_9 ), .A2(n915), .ZN(\U22/Z_9 ) );
  AND2_X1 U367 ( .A1(\U22/DATA1_10 ), .A2(n915), .ZN(\U22/Z_10 ) );
  AND2_X1 U368 ( .A1(\U22/DATA1_11 ), .A2(n915), .ZN(\U22/Z_11 ) );
  AND2_X1 U369 ( .A1(\U22/DATA1_12 ), .A2(n915), .ZN(\U22/Z_12 ) );
  AND2_X1 U370 ( .A1(\U22/DATA1_13 ), .A2(n915), .ZN(\U22/Z_13 ) );
  AND2_X1 U374 ( .A1(\U22/DATA1_14 ), .A2(n915), .ZN(\U22/Z_14 ) );
  AND2_X1 U375 ( .A1(\U22/DATA1_15 ), .A2(n915), .ZN(\U22/Z_15 ) );
  AND2_X1 U376 ( .A1(\U22/DATA1_16 ), .A2(n915), .ZN(\U22/Z_16 ) );
  AND2_X1 U377 ( .A1(\U22/DATA1_17 ), .A2(n915), .ZN(\U22/Z_17 ) );
  AND2_X1 U378 ( .A1(\U22/DATA1_18 ), .A2(n915), .ZN(\U22/Z_18 ) );
  AND2_X1 U383 ( .A1(\U22/DATA1_19 ), .A2(n915), .ZN(\U22/Z_19 ) );
  AND2_X1 U384 ( .A1(\U22/DATA1_20 ), .A2(n915), .ZN(\U22/Z_20 ) );
  AND2_X1 U385 ( .A1(\U22/DATA1_21 ), .A2(n915), .ZN(\U22/Z_21 ) );
  AND2_X1 U386 ( .A1(\U22/DATA1_22 ), .A2(n915), .ZN(\U22/Z_22 ) );
  AND2_X1 U387 ( .A1(\U22/DATA1_23 ), .A2(n915), .ZN(\U22/Z_23 ) );
  AND2_X1 U388 ( .A1(\U22/DATA1_24 ), .A2(n915), .ZN(\U22/Z_24 ) );
  AND2_X1 U389 ( .A1(\U22/DATA1_25 ), .A2(n915), .ZN(\U22/Z_25 ) );
  AND2_X1 U390 ( .A1(\U22/DATA1_26 ), .A2(n915), .ZN(\U22/Z_26 ) );
  AND2_X1 U392 ( .A1(\U22/DATA1_27 ), .A2(n915), .ZN(\U22/Z_27 ) );
  INV_X4 U393 ( .A(divisor[16]), .ZN(n1247) );
  AND2_X1 U394 ( .A1(\U25/DATA1_7 ), .A2(start), .ZN(\U25/Z_7 ) );
  AND2_X1 U395 ( .A1(\U25/DATA1_8 ), .A2(start), .ZN(\U25/Z_8 ) );
  AND2_X1 U396 ( .A1(\U25/DATA1_9 ), .A2(start), .ZN(\U25/Z_9 ) );
  AND2_X1 U397 ( .A1(\U25/DATA1_10 ), .A2(start), .ZN(\U25/Z_10 ) );
  AND2_X1 U398 ( .A1(\U25/DATA1_11 ), .A2(start), .ZN(\U25/Z_11 ) );
  AND2_X1 U399 ( .A1(\U25/DATA1_12 ), .A2(start), .ZN(\U25/Z_12 ) );
  AND2_X1 U400 ( .A1(\U25/DATA1_13 ), .A2(start), .ZN(\U25/Z_13 ) );
  AND2_X1 U401 ( .A1(\U25/DATA1_14 ), .A2(start), .ZN(\U25/Z_14 ) );
  AND2_X1 U403 ( .A1(\U25/DATA1_15 ), .A2(start), .ZN(\U25/Z_15 ) );
  AND2_X1 U404 ( .A1(\U25/DATA1_16 ), .A2(start), .ZN(\U25/Z_16 ) );
  AND2_X1 U405 ( .A1(\U25/DATA1_17 ), .A2(start), .ZN(\U25/Z_17 ) );
  AND2_X1 U406 ( .A1(\U25/DATA1_18 ), .A2(n1131), .ZN(\U25/Z_18 ) );
  AND2_X1 U407 ( .A1(\U25/DATA1_19 ), .A2(start), .ZN(\U25/Z_19 ) );
  AND2_X1 U408 ( .A1(\U25/DATA1_20 ), .A2(n1131), .ZN(\U25/Z_20 ) );
  AND2_X1 U409 ( .A1(\U25/DATA1_21 ), .A2(start), .ZN(\U25/Z_21 ) );
  AND2_X1 U410 ( .A1(\U25/DATA1_22 ), .A2(n1131), .ZN(\U25/Z_22 ) );
  AND2_X1 U411 ( .A1(\U25/DATA1_23 ), .A2(n1131), .ZN(\U25/Z_23 ) );
  AND2_X1 U412 ( .A1(\U25/DATA1_24 ), .A2(n1131), .ZN(\U25/Z_24 ) );
  AND2_X1 U413 ( .A1(\U25/DATA1_25 ), .A2(n1131), .ZN(\U25/Z_25 ) );
  AND2_X1 U414 ( .A1(\U25/DATA1_26 ), .A2(n1131), .ZN(\U25/Z_26 ) );
  AND2_X1 U415 ( .A1(\U25/DATA1_27 ), .A2(n1131), .ZN(\U25/Z_27 ) );
  NAND3_X2 U416 ( .A1(n1240), .A2(n1239), .A3(n1238), .ZN(n1241) );
  NOR4_X2 U417 ( .A1(n1242), .A2(n1241), .A3(n128), .A4(n129), .ZN(n1246) );
  NOR4_X2 U418 ( .A1(n1244), .A2(n1243), .A3(n118), .A4(n119), .ZN(n1245) );
  NAND2_X2 U419 ( .A1(n1246), .A2(n1245), .ZN(n41) );
  AND2_X1 U420 ( .A1(\U5/DATA1_0 ), .A2(n245), .ZN(\U5/Z_0 ) );
  AND2_X1 U421 ( .A1(\U4/DATA1_1 ), .A2(n41), .ZN(\U4/Z_1 ) );
  AND2_X1 U422 ( .A1(\U8/DATA1_0 ), .A2(n383), .ZN(\U8/Z_0 ) );
  AND2_X1 U423 ( .A1(\U5/DATA1_1 ), .A2(n245), .ZN(\U5/Z_1 ) );
  AND2_X1 U424 ( .A1(\U11/DATA1_0 ), .A2(n519), .ZN(\U11/Z_0 ) );
  AND2_X1 U425 ( .A1(\U8/DATA1_1 ), .A2(n383), .ZN(\U8/Z_1 ) );
  AND2_X1 U426 ( .A1(\U14/DATA1_0 ), .A2(n653), .ZN(\U14/Z_0 ) );
  AND2_X1 U427 ( .A1(\U11/DATA1_1 ), .A2(n519), .ZN(\U11/Z_1 ) );
  AND2_X1 U428 ( .A1(\U17/DATA1_0 ), .A2(n1098), .ZN(\U17/Z_0 ) );
  AND2_X1 U429 ( .A1(\U14/DATA1_1 ), .A2(n653), .ZN(\U14/Z_1 ) );
  AND2_X1 U430 ( .A1(\U20/DATA1_0 ), .A2(n915), .ZN(\U20/Z_0 ) );
  AND2_X1 U431 ( .A1(\U17/DATA1_1 ), .A2(n1098), .ZN(\U17/Z_1 ) );
  AND2_X1 U432 ( .A1(\U20/DATA1_1 ), .A2(n915), .ZN(\U20/Z_1 ) );
  NOR2_X2 U433 ( .A1(n1130), .A2(n1116), .ZN(\U21/Z_16 ) );
  NOR2_X2 U434 ( .A1(n1130), .A2(n1117), .ZN(\U21/Z_17 ) );
  NOR2_X2 U435 ( .A1(n1130), .A2(n1115), .ZN(\U21/Z_18 ) );
  NOR2_X2 U436 ( .A1(n1130), .A2(n1118), .ZN(\U21/Z_19 ) );
endmodule


module Output_Result ( clock, reset_n, DataIn, StartIn, Divisor, StartOut, 
        DataOut );
  input [27:0] DataIn;
  input [19:0] Divisor;
  output [7:0] DataOut;
  input clock, reset_n, StartIn;
  output StartOut;


  pipeline_divider divider ( .clock(clock), .reset_n(reset_n), .start(StartIn), 
        .divided(DataIn), .divisor(Divisor), .q(DataOut), .StartOut(StartOut)
         );
endmodule


module Output_Store ( clock, reset_n, StartIn, ResultIn, WriteBus, 
        WriteAddress, WriteEnable, output_base_offset );
  input [7:0] ResultIn;
  output [127:0] WriteBus;
  output [15:0] WriteAddress;
  input clock, reset_n, StartIn, output_base_offset;
  output WriteEnable;
  wire   \U8/DATA1_0 , \U8/DATA1_1 , \U8/DATA1_2 , \U8/DATA1_3 , \U8/DATA1_4 ,
         \U8/DATA1_5 , \U8/DATA1_6 , \U8/DATA1_7 , \U7/Z_0 , \U7/Z_1 ,
         \U7/Z_2 , \U7/Z_3 , \U6/Z_0 , \U5/DATA2_1 , \U5/DATA2_2 ,
         \U5/DATA2_3 , \U5/DATA2_4 , \U4/DATA2_15 , \sub_63/carry[2] ,
         \sub_63/carry[3] , \sub_63/carry[4] , \sub_63/A[0] , \sub_63/A[1] ,
         \sub_63/A[2] , \sub_63/A[3] , \sub_63/A[4] , \add_55/A[0] ,
         \add_55/A[1] , \add_55/A[2] , \add_55/A[3] , \add_55/A[4] ,
         \add_55/A[5] , \add_55/A[6] , \add_55/A[7] , \add_55/A[8] ,
         \add_55/A[9] , \add_55/A[10] , \add_55/A[11] , \add_55/A[12] ,
         \add_55/A[13] , \add_55/A[14] , \add_55/A[15] , n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n136, n153, n163, n164, n165, n168, n169, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n198, n199, n200, n201, n202, n206, n207, n208, n209, n210,
         n211, n212, n213, n215, n216, n217, n218, n220, n221, n222, n223,
         n225, n226, n228, n229, n232, n233, n234, n235, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n255, n256, n257, n258, n259, n261, n263, n264, n265,
         n267, n268, n269, n270, n271, n272, n274, n275, n276, n277, n278,
         n279, n280, n284, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n313, n314, n316, n317, n318, n319,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n333, n334, n336, n337, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719;
  assign \U8/DATA1_0  = ResultIn[0];
  assign \U8/DATA1_1  = ResultIn[1];
  assign \U8/DATA1_2  = ResultIn[2];
  assign \U8/DATA1_3  = ResultIn[3];
  assign \U8/DATA1_4  = ResultIn[4];
  assign \U8/DATA1_5  = ResultIn[5];
  assign \U8/DATA1_6  = ResultIn[6];
  assign \U8/DATA1_7  = ResultIn[7];
  assign \U4/DATA2_15  = output_base_offset;

  XNOR2_X2 \sub_63/U1_A_1  ( .A(\sub_63/A[1] ), .B(\sub_63/A[0] ), .ZN(
        \U5/DATA2_1 ) );
  OR2_X1 \sub_63/U1_B_1  ( .A1(\sub_63/A[1] ), .A2(\sub_63/A[0] ), .ZN(
        \sub_63/carry[2] ) );
  XNOR2_X2 \sub_63/U1_A_2  ( .A(\sub_63/A[2] ), .B(\sub_63/carry[2] ), .ZN(
        \U5/DATA2_2 ) );
  OR2_X1 \sub_63/U1_B_2  ( .A1(\sub_63/A[2] ), .A2(\sub_63/carry[2] ), .ZN(
        \sub_63/carry[3] ) );
  XNOR2_X2 \sub_63/U1_A_3  ( .A(\sub_63/A[3] ), .B(\sub_63/carry[3] ), .ZN(
        \U5/DATA2_3 ) );
  OR2_X1 \sub_63/U1_B_3  ( .A1(\sub_63/A[3] ), .A2(\sub_63/carry[3] ), .ZN(
        \sub_63/carry[4] ) );
  DFFS_X2 \short_count_reg[0]  ( .D(\U7/Z_0 ), .CK(clock), .SN(reset_n), .Q(
        \sub_63/A[0] ), .QN(n66) );
  DFFS_X2 \short_count_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .SN(n528), .Q(
        \sub_63/A[1] ), .QN(n65) );
  DFFS_X2 \short_count_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .SN(n520), .Q(
        \sub_63/A[2] ), .QN(n64) );
  DFFS_X2 \short_count_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .SN(n529), .Q(
        \sub_63/A[3] ), .QN(n63) );
  SDFFR_X2 \short_count_reg[4]  ( .D(1'b0), .SI(n675), .SE(\U5/DATA2_4 ), .CK(
        clock), .RN(n520), .Q(\sub_63/A[4] ), .QN(n499) );
  OAI22_X2 U29 ( .A1(n705), .A2(n493), .B1(n153), .B2(n124), .ZN(n368) );
  OAI22_X2 U30 ( .A1(n705), .A2(n492), .B1(n153), .B2(n123), .ZN(n369) );
  OAI22_X2 U31 ( .A1(n705), .A2(n491), .B1(n153), .B2(n122), .ZN(n370) );
  OAI22_X2 U37 ( .A1(n494), .A2(n169), .B1(n701), .B2(n120), .ZN(n372) );
  NAND2_X2 U41 ( .A1(WriteBus[10]), .A2(n174), .ZN(n175) );
  NAND2_X2 U43 ( .A1(WriteBus[11]), .A2(n174), .ZN(n176) );
  NAND2_X2 U45 ( .A1(WriteBus[12]), .A2(n174), .ZN(n177) );
  NAND2_X2 U47 ( .A1(WriteBus[13]), .A2(n174), .ZN(n178) );
  NAND2_X2 U49 ( .A1(WriteBus[14]), .A2(n174), .ZN(n179) );
  NOR4_X2 U51 ( .A1(n602), .A2(n713), .A3(n181), .A4(n182), .ZN(n180) );
  NAND2_X2 U53 ( .A1(WriteBus[15]), .A2(n183), .ZN(n184) );
  NAND4_X2 U54 ( .A1(n706), .A2(n185), .A3(n696), .A4(n186), .ZN(n183) );
  NAND3_X2 U56 ( .A1(n190), .A2(n191), .A3(n192), .ZN(n187) );
  NAND2_X2 U61 ( .A1(WriteBus[17]), .A2(n196), .ZN(n198) );
  NAND2_X2 U63 ( .A1(WriteBus[18]), .A2(n196), .ZN(n199) );
  NAND2_X2 U65 ( .A1(WriteBus[19]), .A2(n196), .ZN(n200) );
  NAND2_X2 U67 ( .A1(WriteBus[20]), .A2(n196), .ZN(n201) );
  NAND2_X2 U69 ( .A1(WriteBus[21]), .A2(n196), .ZN(n202) );
  NAND2_X2 U73 ( .A1(WriteBus[22]), .A2(n208), .ZN(n209) );
  NAND2_X2 U75 ( .A1(WriteBus[23]), .A2(n208), .ZN(n210) );
  NAND3_X2 U76 ( .A1(n211), .A2(n212), .A3(n672), .ZN(n208) );
  NAND2_X2 U80 ( .A1(WriteBus[25]), .A2(n213), .ZN(n215) );
  NAND2_X2 U82 ( .A1(WriteBus[26]), .A2(n213), .ZN(n216) );
  NAND2_X2 U84 ( .A1(WriteBus[27]), .A2(n213), .ZN(n217) );
  NAND2_X2 U86 ( .A1(WriteBus[28]), .A2(n213), .ZN(n218) );
  OAI22_X2 U89 ( .A1(n704), .A2(n493), .B1(n220), .B2(n119), .ZN(n392) );
  OAI22_X2 U90 ( .A1(n704), .A2(n492), .B1(n220), .B2(n118), .ZN(n393) );
  OAI22_X2 U91 ( .A1(n704), .A2(n491), .B1(n220), .B2(n117), .ZN(n394) );
  NAND2_X2 U92 ( .A1(n515), .A2(n221), .ZN(n220) );
  NAND4_X2 U93 ( .A1(n717), .A2(n670), .A3(n164), .A4(n222), .ZN(n221) );
  OAI22_X2 U95 ( .A1(n703), .A2(n494), .B1(n223), .B2(n115), .ZN(n396) );
  OAI22_X2 U96 ( .A1(n703), .A2(n497), .B1(n223), .B2(n114), .ZN(n397) );
  OAI22_X2 U97 ( .A1(n703), .A2(n495), .B1(n223), .B2(n113), .ZN(n398) );
  OAI22_X2 U98 ( .A1(n703), .A2(n496), .B1(n223), .B2(n112), .ZN(n399) );
  OAI22_X2 U99 ( .A1(n703), .A2(n493), .B1(n223), .B2(n111), .ZN(n400) );
  OAI22_X2 U100 ( .A1(n703), .A2(n492), .B1(n223), .B2(n110), .ZN(n401) );
  OAI22_X2 U101 ( .A1(n703), .A2(n491), .B1(n223), .B2(n109), .ZN(n402) );
  NAND2_X2 U107 ( .A1(WriteBus[41]), .A2(n226), .ZN(n228) );
  OAI22_X2 U110 ( .A1(n497), .A2(n232), .B1(n700), .B2(n108), .ZN(n405) );
  OAI22_X2 U111 ( .A1(n495), .A2(n232), .B1(n700), .B2(n107), .ZN(n406) );
  OAI22_X2 U112 ( .A1(n496), .A2(n232), .B1(n700), .B2(n106), .ZN(n407) );
  OAI22_X2 U113 ( .A1(n493), .A2(n232), .B1(n700), .B2(n105), .ZN(n408) );
  OAI22_X2 U114 ( .A1(n492), .A2(n232), .B1(n700), .B2(n104), .ZN(n409) );
  OAI22_X2 U115 ( .A1(n491), .A2(n232), .B1(n700), .B2(n103), .ZN(n410) );
  NAND2_X2 U116 ( .A1(n673), .A2(n233), .ZN(n232) );
  NAND2_X2 U123 ( .A1(WriteBus[49]), .A2(n239), .ZN(n240) );
  NAND2_X2 U125 ( .A1(WriteBus[50]), .A2(n239), .ZN(n241) );
  NAND2_X2 U127 ( .A1(WriteBus[51]), .A2(n239), .ZN(n242) );
  NAND2_X2 U129 ( .A1(WriteBus[52]), .A2(n239), .ZN(n243) );
  NAND2_X2 U131 ( .A1(WriteBus[53]), .A2(n239), .ZN(n244) );
  NAND2_X2 U133 ( .A1(WriteBus[54]), .A2(n239), .ZN(n245) );
  NOR3_X2 U135 ( .A1(n248), .A2(n677), .A3(n173), .ZN(n246) );
  NAND2_X2 U137 ( .A1(WriteBus[55]), .A2(n249), .ZN(n250) );
  NAND3_X2 U138 ( .A1(n251), .A2(n252), .A3(n247), .ZN(n249) );
  NAND2_X2 U143 ( .A1(WriteBus[57]), .A2(n253), .ZN(n255) );
  NAND2_X2 U145 ( .A1(WriteBus[58]), .A2(n253), .ZN(n256) );
  NAND2_X2 U147 ( .A1(WriteBus[59]), .A2(n253), .ZN(n257) );
  NAND2_X2 U149 ( .A1(WriteBus[60]), .A2(n253), .ZN(n258) );
  NAND2_X2 U151 ( .A1(WriteBus[61]), .A2(n253), .ZN(n259) );
  OAI22_X2 U155 ( .A1(n492), .A2(n265), .B1(n698), .B2(n101), .ZN(n425) );
  OAI22_X2 U156 ( .A1(n491), .A2(n265), .B1(n698), .B2(n100), .ZN(n426) );
  NAND3_X2 U157 ( .A1(n671), .A2(n185), .A3(n498), .ZN(n265) );
  OAI22_X2 U159 ( .A1(n494), .A2(n267), .B1(n697), .B2(n98), .ZN(n428) );
  OAI22_X2 U160 ( .A1(n497), .A2(n267), .B1(n697), .B2(n97), .ZN(n429) );
  OAI22_X2 U161 ( .A1(n495), .A2(n267), .B1(n697), .B2(n96), .ZN(n430) );
  OAI22_X2 U168 ( .A1(n496), .A2(n268), .B1(n702), .B2(n95), .ZN(n431) );
  NAND3_X2 U169 ( .A1(n252), .A2(n195), .A3(n671), .ZN(n268) );
  OAI22_X2 U170 ( .A1(n710), .A2(n493), .B1(n270), .B2(n94), .ZN(n432) );
  OAI22_X2 U171 ( .A1(n710), .A2(n492), .B1(n270), .B2(n93), .ZN(n433) );
  OAI22_X2 U172 ( .A1(n710), .A2(n491), .B1(n270), .B2(n92), .ZN(n434) );
  OAI22_X2 U175 ( .A1(n709), .A2(n494), .B1(n272), .B2(n90), .ZN(n436) );
  OAI22_X2 U176 ( .A1(n709), .A2(n497), .B1(n272), .B2(n89), .ZN(n437) );
  NAND2_X2 U180 ( .A1(WriteBus[75]), .A2(n275), .ZN(n276) );
  NAND2_X2 U182 ( .A1(WriteBus[76]), .A2(n275), .ZN(n277) );
  NAND2_X2 U184 ( .A1(WriteBus[77]), .A2(n275), .ZN(n278) );
  NAND2_X2 U186 ( .A1(WriteBus[78]), .A2(n275), .ZN(n279) );
  NAND2_X2 U188 ( .A1(WriteBus[79]), .A2(n275), .ZN(n280) );
  OAI22_X2 U192 ( .A1(n494), .A2(n284), .B1(n699), .B2(n87), .ZN(n444) );
  NAND3_X2 U193 ( .A1(n238), .A2(n211), .A3(n673), .ZN(n284) );
  NAND2_X2 U196 ( .A1(WriteBus[82]), .A2(n287), .ZN(n288) );
  NAND2_X2 U198 ( .A1(WriteBus[83]), .A2(n287), .ZN(n289) );
  NAND2_X2 U200 ( .A1(WriteBus[84]), .A2(n287), .ZN(n290) );
  NAND2_X2 U202 ( .A1(WriteBus[85]), .A2(n287), .ZN(n291) );
  NAND2_X2 U204 ( .A1(WriteBus[86]), .A2(n287), .ZN(n292) );
  NAND2_X2 U206 ( .A1(WriteBus[87]), .A2(n287), .ZN(n293) );
  NAND2_X2 U209 ( .A1(n163), .A2(n168), .ZN(n296) );
  NAND3_X2 U210 ( .A1(n264), .A2(n297), .A3(n274), .ZN(n295) );
  NAND2_X2 U218 ( .A1(WriteBus[89]), .A2(n301), .ZN(n302) );
  NAND2_X2 U220 ( .A1(WriteBus[90]), .A2(n301), .ZN(n303) );
  NAND2_X2 U222 ( .A1(WriteBus[91]), .A2(n301), .ZN(n304) );
  NAND2_X2 U224 ( .A1(WriteBus[92]), .A2(n301), .ZN(n305) );
  NAND2_X2 U226 ( .A1(WriteBus[93]), .A2(n301), .ZN(n306) );
  NAND2_X2 U228 ( .A1(WriteBus[94]), .A2(n301), .ZN(n307) );
  NAND2_X2 U232 ( .A1(WriteBus[95]), .A2(n310), .ZN(n311) );
  NAND2_X2 U238 ( .A1(WriteBus[97]), .A2(n314), .ZN(n316) );
  NAND2_X2 U240 ( .A1(WriteBus[98]), .A2(n314), .ZN(n317) );
  NAND2_X2 U242 ( .A1(WriteBus[99]), .A2(n314), .ZN(n318) );
  NAND2_X2 U244 ( .A1(WriteBus[100]), .A2(n314), .ZN(n319) );
  NAND2_X2 U247 ( .A1(WriteBus[101]), .A2(n321), .ZN(n322) );
  NAND4_X2 U248 ( .A1(n247), .A2(n323), .A3(n324), .A4(n252), .ZN(n321) );
  NOR2_X2 U249 ( .A1(n286), .A2(n300), .ZN(n324) );
  NAND2_X2 U252 ( .A1(n325), .A2(n190), .ZN(n234) );
  OAI22_X2 U253 ( .A1(n716), .A2(n492), .B1(n326), .B2(n86), .ZN(n465) );
  OAI22_X2 U254 ( .A1(n716), .A2(n491), .B1(n326), .B2(n85), .ZN(n466) );
  OAI22_X2 U257 ( .A1(n715), .A2(n494), .B1(n328), .B2(n83), .ZN(n468) );
  OAI22_X2 U258 ( .A1(n715), .A2(n497), .B1(n328), .B2(n82), .ZN(n469) );
  OAI22_X2 U259 ( .A1(n715), .A2(n495), .B1(n328), .B2(n81), .ZN(n470) );
  OAI22_X2 U262 ( .A1(n496), .A2(n330), .B1(n707), .B2(n80), .ZN(n471) );
  OAI22_X2 U265 ( .A1(n493), .A2(n711), .B1(n333), .B2(n79), .ZN(n472) );
  OAI22_X2 U266 ( .A1(n492), .A2(n711), .B1(n333), .B2(n78), .ZN(n473) );
  OAI22_X2 U267 ( .A1(n491), .A2(n711), .B1(n333), .B2(n77), .ZN(n474) );
  NOR2_X2 U268 ( .A1(n334), .A2(n189), .ZN(n333) );
  NAND2_X2 U269 ( .A1(n247), .A2(n712), .ZN(n189) );
  OAI22_X2 U272 ( .A1(n494), .A2(n337), .B1(n708), .B2(n75), .ZN(n476) );
  OAI22_X2 U273 ( .A1(n497), .A2(n337), .B1(n708), .B2(n74), .ZN(n477) );
  NOR2_X2 U278 ( .A1(n676), .A2(n517), .ZN(n336) );
  NOR3_X2 U281 ( .A1(n173), .A2(n600), .A3(n718), .ZN(n339) );
  NAND2_X2 U282 ( .A1(n325), .A2(n168), .ZN(n207) );
  NOR2_X2 U283 ( .A1(n181), .A2(n679), .ZN(n325) );
  NAND2_X2 U285 ( .A1(WriteBus[115]), .A2(n341), .ZN(n342) );
  NAND2_X2 U287 ( .A1(WriteBus[116]), .A2(n341), .ZN(n343) );
  NAND2_X2 U289 ( .A1(WriteBus[117]), .A2(n341), .ZN(n344) );
  NAND2_X2 U291 ( .A1(WriteBus[118]), .A2(n341), .ZN(n345) );
  NAND2_X2 U293 ( .A1(WriteBus[119]), .A2(n341), .ZN(n346) );
  NOR4_X2 U296 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(n309) );
  NOR2_X2 U304 ( .A1(n679), .A2(n681), .ZN(n351) );
  NAND3_X2 U305 ( .A1(n340), .A2(n194), .A3(n163), .ZN(n172) );
  NOR2_X2 U306 ( .A1(n678), .A2(n677), .ZN(n163) );
  OAI22_X2 U308 ( .A1(n494), .A2(n353), .B1(n714), .B2(n73), .ZN(n484) );
  OAI22_X2 U310 ( .A1(n497), .A2(n353), .B1(n714), .B2(n72), .ZN(n485) );
  OAI22_X2 U312 ( .A1(n495), .A2(n353), .B1(n714), .B2(n71), .ZN(n486) );
  OAI22_X2 U314 ( .A1(n496), .A2(n353), .B1(n714), .B2(n70), .ZN(n487) );
  OAI22_X2 U316 ( .A1(n493), .A2(n353), .B1(n714), .B2(n69), .ZN(n488) );
  OAI22_X2 U318 ( .A1(n492), .A2(n353), .B1(n714), .B2(n68), .ZN(n489) );
  OAI22_X2 U320 ( .A1(n491), .A2(n353), .B1(n714), .B2(n67), .ZN(n490) );
  NAND3_X2 U321 ( .A1(n354), .A2(n261), .A3(n668), .ZN(n353) );
  NAND3_X2 U324 ( .A1(n164), .A2(n352), .A3(n717), .ZN(n355) );
  NAND2_X2 U325 ( .A1(n165), .A2(n194), .ZN(n206) );
  NAND3_X2 U326 ( .A1(n65), .A2(n64), .A3(n356), .ZN(n165) );
  NAND2_X2 U327 ( .A1(n357), .A2(n356), .ZN(n352) );
  NAND3_X2 U328 ( .A1(n66), .A2(n63), .A3(n357), .ZN(n340) );
  NAND3_X2 U329 ( .A1(n65), .A2(n63), .A3(n358), .ZN(n235) );
  NAND3_X2 U330 ( .A1(n356), .A2(n65), .A3(\sub_63/A[2] ), .ZN(n225) );
  NAND3_X2 U334 ( .A1(\sub_63/A[1] ), .A2(n63), .A3(n358), .ZN(n222) );
  NAND3_X2 U335 ( .A1(\sub_63/A[1] ), .A2(n356), .A3(\sub_63/A[2] ), .ZN(n297)
         );
  NOR2_X2 U336 ( .A1(n66), .A2(\sub_63/A[3] ), .ZN(n356) );
  NAND3_X2 U339 ( .A1(n190), .A2(n191), .A3(n329), .ZN(n263) );
  NAND3_X2 U340 ( .A1(\sub_63/A[3] ), .A2(\sub_63/A[1] ), .A3(n358), .ZN(n329)
         );
  NAND3_X2 U341 ( .A1(\sub_63/A[0] ), .A2(n64), .A3(n359), .ZN(n191) );
  NAND3_X2 U342 ( .A1(\sub_63/A[3] ), .A2(n66), .A3(n357), .ZN(n190) );
  NOR2_X2 U345 ( .A1(n64), .A2(\sub_63/A[0] ), .ZN(n358) );
  NAND3_X2 U346 ( .A1(\sub_63/A[3] ), .A2(\sub_63/A[0] ), .A3(n357), .ZN(n274)
         );
  NOR2_X2 U347 ( .A1(n65), .A2(\sub_63/A[2] ), .ZN(n357) );
  NAND3_X2 U348 ( .A1(\sub_63/A[2] ), .A2(\sub_63/A[0] ), .A3(n359), .ZN(n192)
         );
  NOR2_X2 U349 ( .A1(n63), .A2(\sub_63/A[1] ), .ZN(n359) );
  NAND2_X2 U351 ( .A1(\sub_63/A[0] ), .A2(n675), .ZN(\U7/Z_0 ) );
  NOR2_X2 U353 ( .A1(n517), .A2(n360), .ZN(\U6/Z_0 ) );
  NAND4_X2 U354 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(n194) );
  AND2_X1 U421 ( .A1(n313), .A2(n261), .ZN(n247) );
  OR2_X1 U422 ( .A1(n207), .A2(n681), .ZN(n173) );
  AND2_X1 U423 ( .A1(n168), .A2(n340), .ZN(n164) );
  AND2_X1 U424 ( .A1(n225), .A2(n235), .ZN(n168) );
  OR2_X1 U425 ( .A1(\U5/DATA2_3 ), .A2(n136), .ZN(\U7/Z_3 ) );
  OR2_X1 U426 ( .A1(\U5/DATA2_2 ), .A2(n136), .ZN(\U7/Z_2 ) );
  OR2_X1 U427 ( .A1(\U5/DATA2_1 ), .A2(n136), .ZN(\U7/Z_1 ) );
  DFFR_X2 \WriteBus_reg[81]  ( .D(n444), .CK(clock), .RN(n521), .Q(
        WriteBus[81]), .QN(n87) );
  DFFR_X2 \WriteBus_reg[68]  ( .D(n431), .CK(clock), .RN(n523), .Q(
        WriteBus[68]), .QN(n95) );
  DFFR_X2 \WriteBus_reg[9]  ( .D(n372), .CK(clock), .RN(n528), .Q(WriteBus[9]), 
        .QN(n120) );
  DFFR_X2 \WriteBus_reg[127]  ( .D(n490), .CK(clock), .RN(n519), .Q(
        WriteBus[127]), .QN(n67) );
  DFFR_X2 \WriteBus_reg[126]  ( .D(n489), .CK(clock), .RN(n519), .Q(
        WriteBus[126]), .QN(n68) );
  DFFR_X2 \WriteBus_reg[125]  ( .D(n488), .CK(clock), .RN(n519), .Q(
        WriteBus[125]), .QN(n69) );
  DFFR_X2 \WriteBus_reg[124]  ( .D(n487), .CK(clock), .RN(n519), .Q(
        WriteBus[124]), .QN(n70) );
  DFFR_X2 \WriteBus_reg[123]  ( .D(n486), .CK(clock), .RN(n519), .Q(
        WriteBus[123]), .QN(n71) );
  DFFR_X2 \WriteBus_reg[122]  ( .D(n485), .CK(clock), .RN(n519), .Q(
        WriteBus[122]), .QN(n72) );
  DFFR_X2 \WriteBus_reg[121]  ( .D(n484), .CK(clock), .RN(n519), .Q(
        WriteBus[121]), .QN(n73) );
  DFFR_X2 \WriteBus_reg[114]  ( .D(n477), .CK(clock), .RN(n520), .Q(
        WriteBus[114]), .QN(n74) );
  DFFR_X2 \WriteBus_reg[113]  ( .D(n476), .CK(clock), .RN(n520), .Q(
        WriteBus[113]), .QN(n75) );
  DFFR_X2 \WriteBus_reg[111]  ( .D(n474), .CK(clock), .RN(n520), .Q(
        WriteBus[111]), .QN(n77) );
  DFFR_X2 \WriteBus_reg[110]  ( .D(n473), .CK(clock), .RN(n520), .Q(
        WriteBus[110]), .QN(n78) );
  DFFR_X2 \WriteBus_reg[109]  ( .D(n472), .CK(clock), .RN(n520), .Q(
        WriteBus[109]), .QN(n79) );
  DFFR_X2 \WriteBus_reg[108]  ( .D(n471), .CK(clock), .RN(n520), .Q(
        WriteBus[108]), .QN(n80) );
  DFFR_X2 \WriteBus_reg[107]  ( .D(n470), .CK(clock), .RN(n520), .Q(
        WriteBus[107]), .QN(n81) );
  DFFR_X2 \WriteBus_reg[106]  ( .D(n469), .CK(clock), .RN(n520), .Q(
        WriteBus[106]), .QN(n82) );
  DFFR_X2 \WriteBus_reg[105]  ( .D(n468), .CK(clock), .RN(n523), .Q(
        WriteBus[105]), .QN(n83) );
  DFFR_X2 \WriteBus_reg[103]  ( .D(n466), .CK(clock), .RN(n522), .Q(
        WriteBus[103]), .QN(n85) );
  DFFR_X2 \WriteBus_reg[102]  ( .D(n465), .CK(clock), .RN(n528), .Q(
        WriteBus[102]), .QN(n86) );
  DFFR_X2 \WriteBus_reg[74]  ( .D(n437), .CK(clock), .RN(n522), .Q(
        WriteBus[74]), .QN(n89) );
  DFFR_X2 \WriteBus_reg[73]  ( .D(n436), .CK(clock), .RN(n522), .Q(
        WriteBus[73]), .QN(n90) );
  DFFR_X2 \WriteBus_reg[71]  ( .D(n434), .CK(clock), .RN(n522), .Q(
        WriteBus[71]), .QN(n92) );
  DFFR_X2 \WriteBus_reg[70]  ( .D(n433), .CK(clock), .RN(n522), .Q(
        WriteBus[70]), .QN(n93) );
  DFFR_X2 \WriteBus_reg[69]  ( .D(n432), .CK(clock), .RN(n522), .Q(
        WriteBus[69]), .QN(n94) );
  DFFR_X2 \WriteBus_reg[67]  ( .D(n430), .CK(clock), .RN(n523), .Q(
        WriteBus[67]), .QN(n96) );
  DFFR_X2 \WriteBus_reg[66]  ( .D(n429), .CK(clock), .RN(n523), .Q(
        WriteBus[66]), .QN(n97) );
  DFFR_X2 \WriteBus_reg[65]  ( .D(n428), .CK(clock), .RN(n523), .Q(
        WriteBus[65]), .QN(n98) );
  DFFR_X2 \WriteBus_reg[63]  ( .D(n426), .CK(clock), .RN(n523), .Q(
        WriteBus[63]), .QN(n100) );
  DFFR_X2 \WriteBus_reg[62]  ( .D(n425), .CK(clock), .RN(n523), .Q(
        WriteBus[62]), .QN(n101) );
  DFFR_X2 \WriteBus_reg[47]  ( .D(n410), .CK(clock), .RN(n524), .Q(
        WriteBus[47]), .QN(n103) );
  DFFR_X2 \WriteBus_reg[46]  ( .D(n409), .CK(clock), .RN(n524), .Q(
        WriteBus[46]), .QN(n104) );
  DFFR_X2 \WriteBus_reg[45]  ( .D(n408), .CK(clock), .RN(n525), .Q(
        WriteBus[45]), .QN(n105) );
  DFFR_X2 \WriteBus_reg[44]  ( .D(n407), .CK(clock), .RN(n525), .Q(
        WriteBus[44]), .QN(n106) );
  DFFR_X2 \WriteBus_reg[43]  ( .D(n406), .CK(clock), .RN(n525), .Q(
        WriteBus[43]), .QN(n107) );
  DFFR_X2 \WriteBus_reg[42]  ( .D(n405), .CK(clock), .RN(n525), .Q(
        WriteBus[42]), .QN(n108) );
  DFFR_X2 \WriteBus_reg[39]  ( .D(n402), .CK(clock), .RN(n525), .Q(
        WriteBus[39]), .QN(n109) );
  DFFR_X2 \WriteBus_reg[38]  ( .D(n401), .CK(clock), .RN(n525), .Q(
        WriteBus[38]), .QN(n110) );
  DFFR_X2 \WriteBus_reg[37]  ( .D(n400), .CK(clock), .RN(n525), .Q(
        WriteBus[37]), .QN(n111) );
  DFFR_X2 \WriteBus_reg[36]  ( .D(n399), .CK(clock), .RN(n525), .Q(
        WriteBus[36]), .QN(n112) );
  DFFR_X2 \WriteBus_reg[35]  ( .D(n398), .CK(clock), .RN(n525), .Q(
        WriteBus[35]), .QN(n113) );
  DFFR_X2 \WriteBus_reg[34]  ( .D(n397), .CK(clock), .RN(n525), .Q(
        WriteBus[34]), .QN(n114) );
  DFFR_X2 \WriteBus_reg[33]  ( .D(n396), .CK(clock), .RN(n526), .Q(
        WriteBus[33]), .QN(n115) );
  DFFR_X2 \WriteBus_reg[31]  ( .D(n394), .CK(clock), .RN(n526), .Q(
        WriteBus[31]), .QN(n117) );
  DFFR_X2 \WriteBus_reg[30]  ( .D(n393), .CK(clock), .RN(n526), .Q(
        WriteBus[30]), .QN(n118) );
  DFFR_X2 \WriteBus_reg[29]  ( .D(n392), .CK(clock), .RN(n526), .Q(
        WriteBus[29]), .QN(n119) );
  DFFR_X2 \WriteBus_reg[7]  ( .D(n370), .CK(clock), .RN(n528), .Q(WriteBus[7]), 
        .QN(n122) );
  DFFR_X2 \WriteBus_reg[6]  ( .D(n369), .CK(clock), .RN(n528), .Q(WriteBus[6]), 
        .QN(n123) );
  DFFR_X2 \WriteBus_reg[5]  ( .D(n368), .CK(clock), .RN(n527), .Q(WriteBus[5]), 
        .QN(n124) );
  DFFR_X2 \WriteBus_reg[4]  ( .D(n367), .CK(clock), .RN(n528), .Q(WriteBus[4]), 
        .QN(n125) );
  DFFR_X2 \WriteBus_reg[3]  ( .D(n366), .CK(clock), .RN(n528), .Q(WriteBus[3]), 
        .QN(n126) );
  DFFR_X2 \WriteBus_reg[2]  ( .D(n365), .CK(clock), .RN(n528), .Q(WriteBus[2]), 
        .QN(n127) );
  DFFR_X2 \WriteBus_reg[1]  ( .D(n364), .CK(clock), .RN(n528), .Q(WriteBus[1]), 
        .QN(n128) );
  DFFR_X2 \WriteBus_reg[64]  ( .D(n427), .CK(clock), .RN(n523), .Q(
        WriteBus[64]), .QN(n99) );
  DFFR_X2 \WriteBus_reg[112]  ( .D(n475), .CK(clock), .RN(n520), .Q(
        WriteBus[112]), .QN(n76) );
  DFFR_X2 \WriteBus_reg[0]  ( .D(n363), .CK(clock), .RN(n528), .Q(WriteBus[0]), 
        .QN(n129) );
  DFFR_X2 \WriteBus_reg[8]  ( .D(n371), .CK(clock), .RN(n528), .Q(WriteBus[8]), 
        .QN(n121) );
  DFFR_X2 \WriteBus_reg[32]  ( .D(n395), .CK(clock), .RN(n526), .Q(
        WriteBus[32]), .QN(n116) );
  DFFR_X2 \WriteBus_reg[72]  ( .D(n435), .CK(clock), .RN(n522), .Q(
        WriteBus[72]), .QN(n91) );
  DFFR_X2 \WriteBus_reg[104]  ( .D(n467), .CK(clock), .RN(n524), .Q(
        WriteBus[104]), .QN(n84) );
  DFFR_X2 \WriteBus_reg[80]  ( .D(n443), .CK(clock), .RN(n522), .Q(
        WriteBus[80]), .QN(n88) );
  DFF_X2 \WriteAddress_reg[15]  ( .D(\add_55/A[15] ), .CK(clock), .Q(
        WriteAddress[15]) );
  DFF_X2 \WriteAddress_reg[14]  ( .D(\add_55/A[14] ), .CK(clock), .Q(
        WriteAddress[14]) );
  DFF_X2 \WriteAddress_reg[13]  ( .D(\add_55/A[13] ), .CK(clock), .Q(
        WriteAddress[13]) );
  DFF_X2 \WriteAddress_reg[12]  ( .D(\add_55/A[12] ), .CK(clock), .Q(
        WriteAddress[12]) );
  DFF_X2 \WriteAddress_reg[11]  ( .D(\add_55/A[11] ), .CK(clock), .Q(
        WriteAddress[11]) );
  DFF_X2 \WriteAddress_reg[10]  ( .D(\add_55/A[10] ), .CK(clock), .Q(
        WriteAddress[10]) );
  DFF_X2 \WriteAddress_reg[9]  ( .D(\add_55/A[9] ), .CK(clock), .Q(
        WriteAddress[9]) );
  DFF_X2 \WriteAddress_reg[8]  ( .D(\add_55/A[8] ), .CK(clock), .Q(
        WriteAddress[8]) );
  DFF_X2 \WriteAddress_reg[7]  ( .D(\add_55/A[7] ), .CK(clock), .Q(
        WriteAddress[7]) );
  DFF_X2 \WriteAddress_reg[6]  ( .D(\add_55/A[6] ), .CK(clock), .Q(
        WriteAddress[6]) );
  DFF_X2 \WriteAddress_reg[5]  ( .D(\add_55/A[5] ), .CK(clock), .Q(
        WriteAddress[5]) );
  DFF_X2 \WriteAddress_reg[4]  ( .D(\add_55/A[4] ), .CK(clock), .Q(
        WriteAddress[4]) );
  DFF_X2 \WriteAddress_reg[3]  ( .D(\add_55/A[3] ), .CK(clock), .Q(
        WriteAddress[3]) );
  DFF_X2 \WriteAddress_reg[2]  ( .D(\add_55/A[2] ), .CK(clock), .Q(
        WriteAddress[2]) );
  DFF_X2 \WriteAddress_reg[1]  ( .D(\add_55/A[1] ), .CK(clock), .Q(
        WriteAddress[1]) );
  DFF_X2 \WriteAddress_reg[0]  ( .D(\add_55/A[0] ), .CK(clock), .Q(
        WriteAddress[0]) );
  DFFR_X2 \WriteBus_reg[48]  ( .D(n411), .CK(clock), .RN(n524), .Q(
        WriteBus[48]), .QN(n102) );
  DFFR_X2 \next_WriteAddress_reg[0]  ( .D(n362), .CK(clock), .RN(n528), .Q(
        \add_55/A[0] ), .QN(n532) );
  DFFR_X2 \next_WriteAddress_reg[15]  ( .D(n361), .CK(clock), .RN(n519), .Q(
        \add_55/A[15] ), .QN(n595) );
  DFFR_X2 \next_WriteAddress_reg[11]  ( .D(n692), .CK(clock), .RN(n529), .Q(
        \add_55/A[11] ) );
  DFFR_X2 \next_WriteAddress_reg[9]  ( .D(n690), .CK(clock), .RN(n529), .Q(
        \add_55/A[9] ) );
  DFFR_X2 \next_WriteAddress_reg[7]  ( .D(n688), .CK(clock), .RN(n529), .Q(
        \add_55/A[7] ) );
  DFFR_X2 \next_WriteAddress_reg[5]  ( .D(n686), .CK(clock), .RN(n529), .Q(
        \add_55/A[5] ) );
  DFFR_X2 \next_WriteAddress_reg[3]  ( .D(n684), .CK(clock), .RN(n529), .Q(
        \add_55/A[3] ) );
  DFFR_X2 \next_WriteAddress_reg[1]  ( .D(n682), .CK(clock), .RN(n529), .Q(
        \add_55/A[1] ) );
  DFFR_X2 \next_WriteAddress_reg[12]  ( .D(n693), .CK(clock), .RN(n529), .Q(
        \add_55/A[12] ), .QN(n581) );
  DFFR_X2 \next_WriteAddress_reg[10]  ( .D(n691), .CK(clock), .RN(n529), .Q(
        \add_55/A[10] ), .QN(n572) );
  DFFR_X2 \next_WriteAddress_reg[8]  ( .D(n689), .CK(clock), .RN(n529), .Q(
        \add_55/A[8] ), .QN(n563) );
  DFFR_X2 \next_WriteAddress_reg[6]  ( .D(n687), .CK(clock), .RN(n528), .Q(
        \add_55/A[6] ), .QN(n554) );
  DFFR_X2 \next_WriteAddress_reg[4]  ( .D(n685), .CK(clock), .RN(n529), .Q(
        \add_55/A[4] ), .QN(n545) );
  DFFR_X2 \next_WriteAddress_reg[2]  ( .D(n683), .CK(clock), .RN(n529), .Q(
        \add_55/A[2] ), .QN(n537) );
  DFFR_X2 \next_WriteAddress_reg[13]  ( .D(n694), .CK(clock), .RN(n519), .Q(
        \add_55/A[13] ), .QN(n585) );
  DFFR_X2 \next_WriteAddress_reg[14]  ( .D(n695), .CK(clock), .RN(n529), .Q(
        \add_55/A[14] ), .QN(n591) );
  DFFR_X2 WriteEnable_reg ( .D(\U6/Z_0 ), .CK(clock), .RN(n519), .Q(
        WriteEnable) );
  DFFR_X2 \WriteBus_reg[55]  ( .D(n418), .CK(clock), .RN(n524), .Q(
        WriteBus[55]) );
  DFFR_X2 \WriteBus_reg[22]  ( .D(n385), .CK(clock), .RN(n526), .Q(
        WriteBus[22]) );
  DFFR_X2 \WriteBus_reg[23]  ( .D(n386), .CK(clock), .RN(n526), .Q(
        WriteBus[23]) );
  DFFR_X2 \WriteBus_reg[101]  ( .D(n464), .CK(clock), .RN(n521), .Q(
        WriteBus[101]) );
  DFFR_X2 \WriteBus_reg[98]  ( .D(n461), .CK(clock), .RN(n520), .Q(
        WriteBus[98]) );
  DFFR_X2 \WriteBus_reg[100]  ( .D(n463), .CK(clock), .RN(reset_n), .Q(
        WriteBus[100]) );
  DFFR_X2 \WriteBus_reg[99]  ( .D(n462), .CK(clock), .RN(n525), .Q(
        WriteBus[99]) );
  DFFR_X2 \WriteBus_reg[97]  ( .D(n460), .CK(clock), .RN(n524), .Q(
        WriteBus[97]) );
  DFFR_X2 \WriteBus_reg[10]  ( .D(n373), .CK(clock), .RN(n528), .Q(
        WriteBus[10]) );
  DFFR_X2 \WriteBus_reg[12]  ( .D(n375), .CK(clock), .RN(n527), .Q(
        WriteBus[12]) );
  DFFR_X2 \WriteBus_reg[11]  ( .D(n374), .CK(clock), .RN(n527), .Q(
        WriteBus[11]) );
  DFFR_X2 \WriteBus_reg[13]  ( .D(n376), .CK(clock), .RN(n527), .Q(
        WriteBus[13]) );
  DFFR_X2 \WriteBus_reg[14]  ( .D(n377), .CK(clock), .RN(n527), .Q(
        WriteBus[14]) );
  DFFR_X2 \WriteBus_reg[95]  ( .D(n458), .CK(clock), .RN(n529), .Q(
        WriteBus[95]) );
  DFFR_X2 \WriteBus_reg[116]  ( .D(n479), .CK(clock), .RN(n520), .Q(
        WriteBus[116]) );
  DFFR_X2 \WriteBus_reg[115]  ( .D(n478), .CK(clock), .RN(n520), .Q(
        WriteBus[115]) );
  DFFR_X2 \WriteBus_reg[82]  ( .D(n445), .CK(clock), .RN(n521), .Q(
        WriteBus[82]) );
  DFFR_X2 \WriteBus_reg[84]  ( .D(n447), .CK(clock), .RN(n521), .Q(
        WriteBus[84]) );
  DFFR_X2 \WriteBus_reg[83]  ( .D(n446), .CK(clock), .RN(n521), .Q(
        WriteBus[83]) );
  DFFR_X2 \WriteBus_reg[117]  ( .D(n480), .CK(clock), .RN(n520), .Q(
        WriteBus[117]) );
  DFFR_X2 \WriteBus_reg[118]  ( .D(n481), .CK(clock), .RN(n519), .Q(
        WriteBus[118]) );
  DFFR_X2 \WriteBus_reg[119]  ( .D(n482), .CK(clock), .RN(n519), .Q(
        WriteBus[119]) );
  DFFR_X2 \WriteBus_reg[85]  ( .D(n448), .CK(clock), .RN(n521), .Q(
        WriteBus[85]) );
  DFFR_X2 \WriteBus_reg[86]  ( .D(n449), .CK(clock), .RN(n521), .Q(
        WriteBus[86]) );
  DFFR_X2 \WriteBus_reg[87]  ( .D(n450), .CK(clock), .RN(n521), .Q(
        WriteBus[87]) );
  DFFR_X2 \WriteBus_reg[28]  ( .D(n391), .CK(clock), .RN(n526), .Q(
        WriteBus[28]) );
  DFFR_X2 \WriteBus_reg[27]  ( .D(n390), .CK(clock), .RN(n526), .Q(
        WriteBus[27]) );
  DFFR_X2 \WriteBus_reg[26]  ( .D(n389), .CK(clock), .RN(n526), .Q(
        WriteBus[26]) );
  DFFR_X2 \WriteBus_reg[25]  ( .D(n388), .CK(clock), .RN(n526), .Q(
        WriteBus[25]) );
  DFFR_X2 \WriteBus_reg[61]  ( .D(n424), .CK(clock), .RN(n523), .Q(
        WriteBus[61]) );
  DFFR_X2 \WriteBus_reg[60]  ( .D(n423), .CK(clock), .RN(n523), .Q(
        WriteBus[60]) );
  DFFR_X2 \WriteBus_reg[59]  ( .D(n422), .CK(clock), .RN(n523), .Q(
        WriteBus[59]) );
  DFFR_X2 \WriteBus_reg[58]  ( .D(n421), .CK(clock), .RN(n523), .Q(
        WriteBus[58]) );
  DFFR_X2 \WriteBus_reg[57]  ( .D(n420), .CK(clock), .RN(n523), .Q(
        WriteBus[57]) );
  DFFR_X2 \WriteBus_reg[79]  ( .D(n442), .CK(clock), .RN(n522), .Q(
        WriteBus[79]) );
  DFFR_X2 \WriteBus_reg[78]  ( .D(n441), .CK(clock), .RN(n522), .Q(
        WriteBus[78]) );
  DFFR_X2 \WriteBus_reg[77]  ( .D(n440), .CK(clock), .RN(n522), .Q(
        WriteBus[77]) );
  DFFR_X2 \WriteBus_reg[76]  ( .D(n439), .CK(clock), .RN(n522), .Q(
        WriteBus[76]) );
  DFFR_X2 \WriteBus_reg[75]  ( .D(n438), .CK(clock), .RN(n522), .Q(
        WriteBus[75]) );
  DFFR_X2 \WriteBus_reg[15]  ( .D(n378), .CK(clock), .RN(n527), .Q(
        WriteBus[15]) );
  DFFR_X2 \WriteBus_reg[21]  ( .D(n384), .CK(clock), .RN(n527), .Q(
        WriteBus[21]) );
  DFFR_X2 \WriteBus_reg[20]  ( .D(n383), .CK(clock), .RN(n527), .Q(
        WriteBus[20]) );
  DFFR_X2 \WriteBus_reg[19]  ( .D(n382), .CK(clock), .RN(n527), .Q(
        WriteBus[19]) );
  DFFR_X2 \WriteBus_reg[18]  ( .D(n381), .CK(clock), .RN(n527), .Q(
        WriteBus[18]) );
  DFFR_X2 \WriteBus_reg[17]  ( .D(n380), .CK(clock), .RN(n527), .Q(
        WriteBus[17]) );
  DFFR_X2 \WriteBus_reg[41]  ( .D(n404), .CK(clock), .RN(n525), .Q(
        WriteBus[41]) );
  DFFR_X2 \WriteBus_reg[94]  ( .D(n457), .CK(clock), .RN(n526), .Q(
        WriteBus[94]) );
  DFFR_X2 \WriteBus_reg[93]  ( .D(n456), .CK(clock), .RN(n527), .Q(
        WriteBus[93]) );
  DFFR_X2 \WriteBus_reg[92]  ( .D(n455), .CK(clock), .RN(n521), .Q(
        WriteBus[92]) );
  DFFR_X2 \WriteBus_reg[91]  ( .D(n454), .CK(clock), .RN(n521), .Q(
        WriteBus[91]) );
  DFFR_X2 \WriteBus_reg[90]  ( .D(n453), .CK(clock), .RN(n521), .Q(
        WriteBus[90]) );
  DFFR_X2 \WriteBus_reg[89]  ( .D(n452), .CK(clock), .RN(n521), .Q(
        WriteBus[89]) );
  DFFR_X2 \WriteBus_reg[54]  ( .D(n417), .CK(clock), .RN(n524), .Q(
        WriteBus[54]) );
  DFFR_X2 \WriteBus_reg[53]  ( .D(n416), .CK(clock), .RN(n524), .Q(
        WriteBus[53]) );
  DFFR_X2 \WriteBus_reg[52]  ( .D(n415), .CK(clock), .RN(n524), .Q(
        WriteBus[52]) );
  DFFR_X2 \WriteBus_reg[51]  ( .D(n414), .CK(clock), .RN(n524), .Q(
        WriteBus[51]) );
  DFFR_X2 \WriteBus_reg[50]  ( .D(n413), .CK(clock), .RN(n524), .Q(
        WriteBus[50]) );
  DFFR_X2 \WriteBus_reg[49]  ( .D(n412), .CK(clock), .RN(n524), .Q(
        WriteBus[49]) );
  DFFR_X2 \WriteBus_reg[56]  ( .D(n419), .CK(clock), .RN(n524), .Q(
        WriteBus[56]) );
  DFFR_X2 \WriteBus_reg[88]  ( .D(n451), .CK(clock), .RN(n521), .Q(
        WriteBus[88]) );
  DFFR_X2 \WriteBus_reg[16]  ( .D(n379), .CK(clock), .RN(n527), .Q(
        WriteBus[16]) );
  DFFR_X2 \WriteBus_reg[40]  ( .D(n403), .CK(clock), .RN(n525), .Q(
        WriteBus[40]) );
  DFFR_X2 \WriteBus_reg[96]  ( .D(n459), .CK(clock), .RN(reset_n), .Q(
        WriteBus[96]) );
  DFFR_X2 \WriteBus_reg[24]  ( .D(n387), .CK(clock), .RN(n526), .Q(
        WriteBus[24]) );
  DFFR_X2 \WriteBus_reg[120]  ( .D(n483), .CK(clock), .RN(n519), .Q(
        WriteBus[120]) );
  NAND2_X4 U4 ( .A1(\U8/DATA1_0 ), .A2(n516), .ZN(n512) );
  NAND2_X2 U5 ( .A1(\U8/DATA1_0 ), .A2(n516), .ZN(n659) );
  NAND2_X2 U6 ( .A1(\U8/DATA1_7 ), .A2(n516), .ZN(n491) );
  NAND2_X2 U7 ( .A1(\U8/DATA1_6 ), .A2(n516), .ZN(n492) );
  NAND2_X2 U8 ( .A1(\U8/DATA1_5 ), .A2(n516), .ZN(n493) );
  NAND2_X2 U9 ( .A1(\U8/DATA1_1 ), .A2(n516), .ZN(n494) );
  NAND2_X2 U10 ( .A1(\U8/DATA1_3 ), .A2(n516), .ZN(n495) );
  NAND2_X2 U11 ( .A1(\U8/DATA1_4 ), .A2(n516), .ZN(n496) );
  NAND2_X2 U12 ( .A1(\U8/DATA1_2 ), .A2(n516), .ZN(n497) );
  AND3_X4 U13 ( .A1(n212), .A2(n634), .A3(n633), .ZN(n498) );
  NAND2_X1 U14 ( .A1(n664), .A2(n618), .ZN(n500) );
  NAND2_X2 U15 ( .A1(WriteBus[40]), .A2(n226), .ZN(n501) );
  NAND2_X2 U16 ( .A1(n500), .A2(n501), .ZN(n403) );
  OAI22_X1 U17 ( .A1(n705), .A2(n494), .B1(n153), .B2(n128), .ZN(n364) );
  OAI22_X1 U18 ( .A1(n705), .A2(n497), .B1(n153), .B2(n127), .ZN(n365) );
  OAI22_X1 U19 ( .A1(n705), .A2(n495), .B1(n153), .B2(n126), .ZN(n366) );
  OAI22_X1 U20 ( .A1(n705), .A2(n496), .B1(n153), .B2(n125), .ZN(n367) );
  NOR2_X1 U21 ( .A1(n248), .A2(n309), .ZN(n347) );
  NAND2_X1 U22 ( .A1(n313), .A2(n667), .ZN(n650) );
  NOR4_X1 U23 ( .A1(n309), .A2(n602), .A3(n669), .A4(n263), .ZN(n308) );
  NAND2_X1 U24 ( .A1(n664), .A2(n502), .ZN(n503) );
  NAND2_X2 U25 ( .A1(WriteBus[88]), .A2(n511), .ZN(n504) );
  NAND2_X2 U26 ( .A1(n503), .A2(n504), .ZN(n451) );
  INV_X4 U27 ( .A(n511), .ZN(n502) );
  MUX2_X2 U28 ( .A(n664), .B(WriteBus[24]), .S(n213), .Z(n387) );
  MUX2_X2 U32 ( .A(n664), .B(WriteBus[96]), .S(n314), .Z(n459) );
  NAND2_X1 U33 ( .A1(n664), .A2(n505), .ZN(n506) );
  NAND2_X2 U34 ( .A1(WriteBus[56]), .A2(n253), .ZN(n507) );
  NAND2_X2 U35 ( .A1(n506), .A2(n507), .ZN(n419) );
  INV_X4 U36 ( .A(n253), .ZN(n505) );
  NAND2_X1 U38 ( .A1(n664), .A2(n508), .ZN(n509) );
  NAND2_X2 U39 ( .A1(WriteBus[16]), .A2(n196), .ZN(n510) );
  NAND2_X2 U40 ( .A1(n509), .A2(n510), .ZN(n379) );
  INV_X4 U42 ( .A(n196), .ZN(n508) );
  OR4_X1 U44 ( .A1(n647), .A2(n646), .A3(n645), .A4(n665), .ZN(n511) );
  INV_X2 U46 ( .A(n625), .ZN(n411) );
  INV_X2 U48 ( .A(n643), .ZN(n443) );
  INV_X2 U50 ( .A(n654), .ZN(n467) );
  INV_X2 U52 ( .A(n640), .ZN(n435) );
  INV_X2 U55 ( .A(n616), .ZN(n395) );
  INV_X2 U57 ( .A(n611), .ZN(n371) );
  INV_X2 U58 ( .A(n607), .ZN(n363) );
  INV_X2 U59 ( .A(n660), .ZN(n475) );
  INV_X2 U60 ( .A(n636), .ZN(n427) );
  AND4_X4 U62 ( .A1(n672), .A2(n212), .A3(n612), .A4(n633), .ZN(n513) );
  NAND2_X1 U64 ( .A1(n673), .A2(n171), .ZN(n169) );
  NOR3_X1 U66 ( .A1(n719), .A2(n309), .A3(n669), .ZN(n331) );
  INV_X4 U68 ( .A(n530), .ZN(n521) );
  INV_X4 U70 ( .A(n530), .ZN(n524) );
  INV_X4 U71 ( .A(n530), .ZN(n527) );
  INV_X4 U72 ( .A(n530), .ZN(n526) );
  INV_X4 U74 ( .A(n530), .ZN(n523) );
  INV_X4 U77 ( .A(n530), .ZN(n522) );
  INV_X4 U78 ( .A(n530), .ZN(n520) );
  INV_X4 U79 ( .A(n530), .ZN(n529) );
  INV_X4 U81 ( .A(n530), .ZN(n528) );
  INV_X4 U83 ( .A(n530), .ZN(n525) );
  NAND2_X2 U85 ( .A1(n513), .A2(n631), .ZN(n196) );
  NAND2_X1 U87 ( .A1(n668), .A2(n672), .ZN(n275) );
  INV_X4 U88 ( .A(n530), .ZN(n519) );
  INV_X4 U94 ( .A(reset_n), .ZN(n530) );
  OAI21_X2 U102 ( .B1(n718), .B2(n207), .A(n515), .ZN(n211) );
  OAI211_X1 U103 ( .C1(n246), .C2(n517), .A(n238), .B(n247), .ZN(n239) );
  OAI21_X2 U104 ( .B1(n229), .B2(n234), .A(n515), .ZN(n233) );
  AOI21_X2 U105 ( .B1(n515), .B2(n719), .A(n336), .ZN(n313) );
  OAI21_X2 U106 ( .B1(n602), .B2(n327), .A(n515), .ZN(n326) );
  INV_X4 U108 ( .A(n517), .ZN(n516) );
  OAI21_X1 U109 ( .B1(n229), .B2(n617), .A(n515), .ZN(n618) );
  INV_X4 U117 ( .A(n517), .ZN(n515) );
  AND3_X2 U118 ( .A1(n655), .A2(n656), .A3(n313), .ZN(n514) );
  OAI211_X2 U119 ( .C1(n180), .C2(n517), .A(n712), .B(n706), .ZN(n174) );
  NAND2_X1 U120 ( .A1(n360), .A2(n516), .ZN(n136) );
  OAI21_X1 U121 ( .B1(n680), .B2(n271), .A(n515), .ZN(n270) );
  OAI21_X1 U122 ( .B1(n679), .B2(n678), .A(n515), .ZN(n195) );
  OAI21_X1 U124 ( .B1(n678), .B2(n234), .A(n515), .ZN(n323) );
  OAI211_X1 U126 ( .C1(n308), .C2(n517), .A(n261), .B(n668), .ZN(n301) );
  AOI21_X2 U128 ( .B1(n667), .B2(n347), .A(n517), .ZN(n341) );
  NAND4_X1 U130 ( .A1(n261), .A2(n185), .A3(n629), .A4(n252), .ZN(n253) );
  OAI21_X1 U132 ( .B1(n248), .B2(n263), .A(n515), .ZN(n354) );
  AOI211_X1 U134 ( .C1(n515), .C2(n187), .A(n188), .B(n189), .ZN(n186) );
  NAND2_X2 U136 ( .A1(n513), .A2(n614), .ZN(n213) );
  OAI21_X2 U139 ( .B1(n339), .B2(n517), .A(n238), .ZN(n334) );
  INV_X4 U140 ( .A(StartIn), .ZN(n517) );
  NAND4_X1 U141 ( .A1(n674), .A2(n294), .A3(n238), .A4(n269), .ZN(n287) );
  OAI21_X1 U142 ( .B1(n295), .B2(n296), .A(n515), .ZN(n294) );
  OAI21_X1 U144 ( .B1(n517), .B2(n194), .A(n195), .ZN(n193) );
  OAI211_X1 U146 ( .C1(n331), .C2(n517), .A(n261), .B(n666), .ZN(n330) );
  OAI21_X2 U148 ( .B1(n491), .B2(n183), .A(n184), .ZN(n378) );
  OAI21_X2 U150 ( .B1(n494), .B2(n196), .A(n198), .ZN(n380) );
  OAI21_X2 U152 ( .B1(n497), .B2(n196), .A(n199), .ZN(n381) );
  OAI21_X2 U153 ( .B1(n495), .B2(n196), .A(n200), .ZN(n382) );
  OAI21_X2 U154 ( .B1(n496), .B2(n196), .A(n201), .ZN(n383) );
  OAI21_X2 U158 ( .B1(n493), .B2(n196), .A(n202), .ZN(n384) );
  OAI21_X2 U162 ( .B1(n492), .B2(n208), .A(n209), .ZN(n385) );
  OAI21_X2 U163 ( .B1(n491), .B2(n208), .A(n210), .ZN(n386) );
  OAI21_X2 U164 ( .B1(n494), .B2(n213), .A(n215), .ZN(n388) );
  OAI21_X2 U165 ( .B1(n497), .B2(n213), .A(n216), .ZN(n389) );
  OAI21_X2 U166 ( .B1(n495), .B2(n213), .A(n217), .ZN(n390) );
  OAI21_X2 U167 ( .B1(n496), .B2(n213), .A(n218), .ZN(n391) );
  OAI21_X2 U173 ( .B1(n226), .B2(n494), .A(n228), .ZN(n404) );
  OAI21_X2 U174 ( .B1(n494), .B2(n239), .A(n240), .ZN(n412) );
  OAI21_X2 U177 ( .B1(n497), .B2(n239), .A(n241), .ZN(n413) );
  OAI21_X2 U178 ( .B1(n495), .B2(n239), .A(n242), .ZN(n414) );
  OAI21_X2 U179 ( .B1(n496), .B2(n239), .A(n243), .ZN(n415) );
  OAI21_X2 U181 ( .B1(n493), .B2(n239), .A(n244), .ZN(n416) );
  OAI21_X2 U183 ( .B1(n492), .B2(n239), .A(n245), .ZN(n417) );
  OAI21_X2 U185 ( .B1(n495), .B2(n275), .A(n276), .ZN(n438) );
  OAI21_X2 U187 ( .B1(n496), .B2(n275), .A(n277), .ZN(n439) );
  OAI21_X2 U189 ( .B1(n493), .B2(n275), .A(n278), .ZN(n440) );
  OAI21_X2 U190 ( .B1(n492), .B2(n275), .A(n279), .ZN(n441) );
  OAI21_X2 U191 ( .B1(n491), .B2(n275), .A(n280), .ZN(n442) );
  OAI21_X2 U194 ( .B1(n494), .B2(n301), .A(n302), .ZN(n452) );
  OAI21_X2 U195 ( .B1(n497), .B2(n301), .A(n303), .ZN(n453) );
  OAI21_X2 U197 ( .B1(n495), .B2(n301), .A(n304), .ZN(n454) );
  OAI21_X2 U199 ( .B1(n496), .B2(n301), .A(n305), .ZN(n455) );
  OAI21_X2 U201 ( .B1(n493), .B2(n301), .A(n306), .ZN(n456) );
  OAI21_X2 U203 ( .B1(n492), .B2(n301), .A(n307), .ZN(n457) );
  OAI21_X2 U205 ( .B1(n494), .B2(n314), .A(n316), .ZN(n460) );
  OAI21_X2 U207 ( .B1(n497), .B2(n314), .A(n317), .ZN(n461) );
  OAI21_X2 U208 ( .B1(n495), .B2(n314), .A(n318), .ZN(n462) );
  OAI21_X2 U211 ( .B1(n496), .B2(n314), .A(n319), .ZN(n463) );
  OAI21_X2 U212 ( .B1(n341), .B2(n495), .A(n342), .ZN(n478) );
  OAI21_X2 U213 ( .B1(n341), .B2(n496), .A(n343), .ZN(n479) );
  OAI21_X2 U214 ( .B1(n341), .B2(n493), .A(n344), .ZN(n480) );
  OAI21_X2 U215 ( .B1(n341), .B2(n492), .A(n345), .ZN(n481) );
  OAI21_X2 U216 ( .B1(n341), .B2(n491), .A(n346), .ZN(n482) );
  OAI21_X1 U217 ( .B1(n172), .B2(n173), .A(n515), .ZN(n171) );
  OAI21_X2 U219 ( .B1(n497), .B2(n174), .A(n175), .ZN(n373) );
  OAI21_X2 U221 ( .B1(n495), .B2(n174), .A(n176), .ZN(n374) );
  OAI21_X2 U223 ( .B1(n496), .B2(n174), .A(n177), .ZN(n375) );
  OAI21_X2 U225 ( .B1(n493), .B2(n174), .A(n178), .ZN(n376) );
  OAI21_X2 U227 ( .B1(n492), .B2(n174), .A(n179), .ZN(n377) );
  OAI21_X2 U229 ( .B1(n491), .B2(n249), .A(n250), .ZN(n418) );
  OAI21_X1 U230 ( .B1(n234), .B2(n248), .A(n515), .ZN(n251) );
  OAI21_X2 U231 ( .B1(n494), .B2(n253), .A(n255), .ZN(n420) );
  OAI21_X2 U233 ( .B1(n497), .B2(n253), .A(n256), .ZN(n421) );
  OAI21_X2 U234 ( .B1(n495), .B2(n253), .A(n257), .ZN(n422) );
  OAI21_X2 U235 ( .B1(n496), .B2(n253), .A(n258), .ZN(n423) );
  OAI21_X2 U236 ( .B1(n493), .B2(n253), .A(n259), .ZN(n424) );
  OAI21_X2 U237 ( .B1(n497), .B2(n287), .A(n288), .ZN(n445) );
  OAI21_X2 U239 ( .B1(n495), .B2(n287), .A(n289), .ZN(n446) );
  OAI21_X2 U241 ( .B1(n496), .B2(n287), .A(n290), .ZN(n447) );
  OAI21_X2 U243 ( .B1(n493), .B2(n287), .A(n291), .ZN(n448) );
  OAI21_X2 U245 ( .B1(n492), .B2(n287), .A(n292), .ZN(n449) );
  OAI21_X2 U246 ( .B1(n491), .B2(n287), .A(n293), .ZN(n450) );
  OAI21_X2 U250 ( .B1(n310), .B2(n491), .A(n311), .ZN(n458) );
  AOI21_X1 U251 ( .B1(n514), .B2(n667), .A(n517), .ZN(n310) );
  OAI21_X2 U255 ( .B1(n493), .B2(n321), .A(n322), .ZN(n464) );
  OAI21_X2 U256 ( .B1(n532), .B2(n136), .A(n533), .ZN(n362) );
  INV_X1 U260 ( .A(\U4/DATA2_15 ), .ZN(n518) );
  INV_X4 U261 ( .A(n194), .ZN(n531) );
  NAND2_X2 U263 ( .A1(n499), .A2(n531), .ZN(n360) );
  INV_X4 U264 ( .A(n136), .ZN(n675) );
  XOR2_X2 U270 ( .A(n499), .B(\sub_63/carry[4] ), .Z(\U5/DATA2_4 ) );
  NAND2_X2 U271 ( .A1(n136), .A2(n516), .ZN(n590) );
  INV_X4 U274 ( .A(n590), .ZN(n597) );
  NAND2_X2 U275 ( .A1(n597), .A2(n532), .ZN(n533) );
  NOR2_X2 U276 ( .A1(n590), .A2(n532), .ZN(n534) );
  NAND2_X2 U277 ( .A1(n533), .A2(n136), .ZN(n536) );
  MUX2_X2 U279 ( .A(n534), .B(n536), .S(\add_55/A[1] ), .Z(n682) );
  NAND2_X2 U280 ( .A1(\add_55/A[0] ), .A2(n537), .ZN(n535) );
  MUX2_X2 U284 ( .A(n537), .B(n535), .S(\add_55/A[1] ), .Z(n539) );
  INV_X4 U286 ( .A(n536), .ZN(n538) );
  OAI22_X2 U288 ( .A1(n539), .A2(n590), .B1(n538), .B2(n537), .ZN(n683) );
  NAND3_X2 U290 ( .A1(\add_55/A[1] ), .A2(\add_55/A[0] ), .A3(\add_55/A[2] ), 
        .ZN(n542) );
  NOR2_X2 U292 ( .A1(n590), .A2(n542), .ZN(n541) );
  NAND2_X2 U294 ( .A1(n597), .A2(n542), .ZN(n540) );
  NAND2_X2 U295 ( .A1(n540), .A2(n136), .ZN(n544) );
  MUX2_X2 U297 ( .A(n541), .B(n544), .S(\add_55/A[3] ), .Z(n684) );
  INV_X4 U298 ( .A(n542), .ZN(n548) );
  NAND2_X2 U299 ( .A1(n548), .A2(n545), .ZN(n543) );
  MUX2_X2 U300 ( .A(n545), .B(n543), .S(\add_55/A[3] ), .Z(n547) );
  INV_X4 U301 ( .A(n544), .ZN(n546) );
  OAI22_X2 U302 ( .A1(n547), .A2(n590), .B1(n546), .B2(n545), .ZN(n685) );
  NAND3_X2 U303 ( .A1(\add_55/A[4] ), .A2(\add_55/A[3] ), .A3(n548), .ZN(n551)
         );
  NOR2_X2 U307 ( .A1(n590), .A2(n551), .ZN(n550) );
  NAND2_X2 U309 ( .A1(n597), .A2(n551), .ZN(n549) );
  NAND2_X2 U311 ( .A1(n549), .A2(n136), .ZN(n553) );
  MUX2_X2 U313 ( .A(n550), .B(n553), .S(\add_55/A[5] ), .Z(n686) );
  INV_X4 U315 ( .A(n551), .ZN(n557) );
  NAND2_X2 U317 ( .A1(n557), .A2(n554), .ZN(n552) );
  MUX2_X2 U319 ( .A(n554), .B(n552), .S(\add_55/A[5] ), .Z(n556) );
  INV_X4 U322 ( .A(n553), .ZN(n555) );
  OAI22_X2 U323 ( .A1(n556), .A2(n590), .B1(n555), .B2(n554), .ZN(n687) );
  NAND3_X2 U331 ( .A1(\add_55/A[6] ), .A2(\add_55/A[5] ), .A3(n557), .ZN(n560)
         );
  NOR2_X2 U332 ( .A1(n590), .A2(n560), .ZN(n559) );
  NAND2_X2 U333 ( .A1(n597), .A2(n560), .ZN(n558) );
  NAND2_X2 U337 ( .A1(n558), .A2(n136), .ZN(n562) );
  MUX2_X2 U338 ( .A(n559), .B(n562), .S(\add_55/A[7] ), .Z(n688) );
  INV_X4 U343 ( .A(n560), .ZN(n566) );
  NAND2_X2 U344 ( .A1(n566), .A2(n563), .ZN(n561) );
  MUX2_X2 U350 ( .A(n563), .B(n561), .S(\add_55/A[7] ), .Z(n565) );
  INV_X4 U352 ( .A(n562), .ZN(n564) );
  OAI22_X2 U355 ( .A1(n565), .A2(n590), .B1(n564), .B2(n563), .ZN(n689) );
  NAND3_X2 U356 ( .A1(\add_55/A[8] ), .A2(\add_55/A[7] ), .A3(n566), .ZN(n569)
         );
  NOR2_X2 U357 ( .A1(n590), .A2(n569), .ZN(n568) );
  NAND2_X2 U358 ( .A1(n597), .A2(n569), .ZN(n567) );
  NAND2_X2 U359 ( .A1(n567), .A2(n136), .ZN(n571) );
  MUX2_X2 U360 ( .A(n568), .B(n571), .S(\add_55/A[9] ), .Z(n690) );
  INV_X4 U361 ( .A(n569), .ZN(n575) );
  NAND2_X2 U362 ( .A1(n575), .A2(n572), .ZN(n570) );
  MUX2_X2 U363 ( .A(n572), .B(n570), .S(\add_55/A[9] ), .Z(n574) );
  INV_X4 U364 ( .A(n571), .ZN(n573) );
  OAI22_X2 U365 ( .A1(n574), .A2(n590), .B1(n573), .B2(n572), .ZN(n691) );
  NAND3_X2 U366 ( .A1(\add_55/A[10] ), .A2(\add_55/A[9] ), .A3(n575), .ZN(n578) );
  NOR2_X2 U367 ( .A1(n590), .A2(n578), .ZN(n577) );
  NAND2_X2 U368 ( .A1(n597), .A2(n578), .ZN(n576) );
  NAND2_X2 U369 ( .A1(n576), .A2(n136), .ZN(n580) );
  MUX2_X2 U370 ( .A(n577), .B(n580), .S(\add_55/A[11] ), .Z(n692) );
  INV_X4 U371 ( .A(n578), .ZN(n584) );
  NAND2_X2 U372 ( .A1(n584), .A2(n581), .ZN(n579) );
  MUX2_X2 U373 ( .A(n581), .B(n579), .S(\add_55/A[11] ), .Z(n583) );
  INV_X4 U374 ( .A(n580), .ZN(n582) );
  OAI22_X2 U375 ( .A1(n583), .A2(n590), .B1(n582), .B2(n581), .ZN(n693) );
  NAND3_X2 U376 ( .A1(\add_55/A[11] ), .A2(\add_55/A[12] ), .A3(n584), .ZN(
        n587) );
  XOR2_X2 U377 ( .A(n587), .B(\add_55/A[13] ), .Z(n586) );
  OAI22_X2 U378 ( .A1(n590), .A2(n586), .B1(n136), .B2(n585), .ZN(n694) );
  INV_X4 U379 ( .A(n587), .ZN(n588) );
  NAND2_X2 U380 ( .A1(\add_55/A[13] ), .A2(n588), .ZN(n594) );
  XOR2_X2 U381 ( .A(n594), .B(\add_55/A[14] ), .Z(n589) );
  OAI22_X2 U382 ( .A1(n590), .A2(n589), .B1(n136), .B2(n591), .ZN(n695) );
  NOR2_X2 U383 ( .A1(n591), .A2(n594), .ZN(n592) );
  NOR2_X2 U384 ( .A1(n517), .A2(n592), .ZN(n593) );
  NOR2_X2 U385 ( .A1(n675), .A2(n593), .ZN(n599) );
  INV_X4 U386 ( .A(n594), .ZN(n596) );
  NAND4_X2 U387 ( .A1(\add_55/A[14] ), .A2(n597), .A3(n596), .A4(n595), .ZN(
        n598) );
  OAI221_X2 U388 ( .B1(n595), .B2(n599), .C1(n515), .C2(n518), .A(n598), .ZN(
        n361) );
  INV_X4 U389 ( .A(n274), .ZN(n600) );
  NAND2_X2 U390 ( .A1(n516), .A2(n600), .ZN(n706) );
  INV_X4 U391 ( .A(n191), .ZN(n680) );
  NAND2_X2 U392 ( .A1(n515), .A2(n680), .ZN(n269) );
  NAND3_X2 U393 ( .A1(n64), .A2(n66), .A3(n359), .ZN(n264) );
  INV_X4 U394 ( .A(n264), .ZN(n601) );
  NAND2_X2 U395 ( .A1(n601), .A2(n516), .ZN(n185) );
  INV_X4 U396 ( .A(n192), .ZN(n602) );
  NAND2_X2 U397 ( .A1(n515), .A2(n602), .ZN(n656) );
  INV_X4 U398 ( .A(n189), .ZN(n603) );
  NAND2_X2 U399 ( .A1(n656), .A2(n603), .ZN(n645) );
  INV_X4 U400 ( .A(n645), .ZN(n674) );
  NAND2_X2 U401 ( .A1(n674), .A2(n706), .ZN(n641) );
  INV_X4 U402 ( .A(n641), .ZN(n673) );
  INV_X4 U403 ( .A(n190), .ZN(n681) );
  NAND2_X2 U404 ( .A1(n515), .A2(n681), .ZN(n644) );
  NAND2_X2 U405 ( .A1(n673), .A2(n644), .ZN(n604) );
  INV_X4 U406 ( .A(n604), .ZN(n672) );
  NAND2_X2 U407 ( .A1(n672), .A2(n269), .ZN(n605) );
  INV_X4 U408 ( .A(n605), .ZN(n671) );
  INV_X4 U409 ( .A(n297), .ZN(n679) );
  NAND2_X2 U410 ( .A1(n515), .A2(n679), .ZN(n635) );
  NAND3_X2 U411 ( .A1(n671), .A2(n185), .A3(n635), .ZN(n617) );
  INV_X4 U412 ( .A(n617), .ZN(n670) );
  NAND4_X2 U413 ( .A1(n165), .A2(n163), .A3(n164), .A4(n670), .ZN(n606) );
  NAND2_X2 U414 ( .A1(n606), .A2(n516), .ZN(n153) );
  INV_X4 U415 ( .A(n153), .ZN(n705) );
  MUX2_X2 U416 ( .A(n512), .B(n129), .S(n705), .Z(n607) );
  INV_X4 U417 ( .A(n168), .ZN(n608) );
  NOR3_X2 U418 ( .A1(n172), .A2(n617), .A3(n608), .ZN(n609) );
  NOR2_X2 U419 ( .A1(n517), .A2(n609), .ZN(n610) );
  MUX2_X2 U420 ( .A(n512), .B(n121), .S(n610), .Z(n611) );
  NAND2_X2 U428 ( .A1(n206), .A2(n516), .ZN(n212) );
  NAND2_X2 U429 ( .A1(n207), .A2(n516), .ZN(n612) );
  INV_X4 U430 ( .A(n222), .ZN(n678) );
  NAND2_X2 U431 ( .A1(n516), .A2(n678), .ZN(n633) );
  INV_X4 U432 ( .A(n352), .ZN(n677) );
  NAND2_X2 U433 ( .A1(n516), .A2(n677), .ZN(n631) );
  INV_X4 U434 ( .A(n659), .ZN(n664) );
  INV_X4 U435 ( .A(n340), .ZN(n613) );
  NAND2_X2 U436 ( .A1(n516), .A2(n613), .ZN(n614) );
  INV_X4 U437 ( .A(n172), .ZN(n637) );
  NAND4_X2 U438 ( .A1(n225), .A2(n165), .A3(n670), .A4(n637), .ZN(n615) );
  NAND2_X2 U439 ( .A1(n615), .A2(n516), .ZN(n223) );
  INV_X4 U440 ( .A(n223), .ZN(n703) );
  MUX2_X2 U441 ( .A(n512), .B(n116), .S(n703), .Z(n616) );
  NAND3_X2 U442 ( .A1(n235), .A2(n165), .A3(n637), .ZN(n229) );
  INV_X4 U443 ( .A(n618), .ZN(n226) );
  NAND2_X2 U444 ( .A1(n340), .A2(n717), .ZN(n619) );
  NAND2_X2 U445 ( .A1(n619), .A2(n516), .ZN(n238) );
  INV_X4 U446 ( .A(n631), .ZN(n623) );
  INV_X4 U447 ( .A(n173), .ZN(n620) );
  NOR2_X2 U448 ( .A1(n517), .A2(n620), .ZN(n622) );
  INV_X4 U449 ( .A(n238), .ZN(n621) );
  NOR4_X2 U450 ( .A1(n623), .A2(n622), .A3(n621), .A4(n641), .ZN(n624) );
  MUX2_X2 U451 ( .A(n102), .B(n512), .S(n624), .Z(n625) );
  NAND2_X2 U452 ( .A1(\sub_63/A[4] ), .A2(n516), .ZN(n261) );
  NAND2_X2 U453 ( .A1(n355), .A2(n516), .ZN(n252) );
  NAND2_X2 U454 ( .A1(n358), .A2(n359), .ZN(n655) );
  NAND3_X2 U455 ( .A1(n192), .A2(n274), .A3(n655), .ZN(n248) );
  INV_X4 U456 ( .A(n309), .ZN(n676) );
  INV_X4 U457 ( .A(n248), .ZN(n627) );
  INV_X4 U458 ( .A(n263), .ZN(n626) );
  NAND4_X2 U459 ( .A1(n222), .A2(n676), .A3(n627), .A4(n626), .ZN(n628) );
  NAND2_X2 U460 ( .A1(n628), .A2(n516), .ZN(n629) );
  INV_X4 U461 ( .A(n164), .ZN(n630) );
  NAND2_X2 U462 ( .A1(n516), .A2(n630), .ZN(n632) );
  NAND2_X2 U463 ( .A1(n632), .A2(n631), .ZN(n188) );
  INV_X4 U464 ( .A(n188), .ZN(n634) );
  NAND3_X2 U465 ( .A1(n498), .A2(n671), .A3(n635), .ZN(n267) );
  INV_X4 U466 ( .A(n267), .ZN(n697) );
  MUX2_X2 U467 ( .A(n99), .B(n512), .S(n697), .Z(n636) );
  NAND4_X2 U468 ( .A1(n351), .A2(n168), .A3(n261), .A4(n637), .ZN(n182) );
  INV_X4 U469 ( .A(n182), .ZN(n649) );
  NAND4_X2 U470 ( .A1(n274), .A2(n165), .A3(n514), .A4(n649), .ZN(n271) );
  INV_X4 U471 ( .A(n271), .ZN(n638) );
  NAND2_X2 U472 ( .A1(n264), .A2(n638), .ZN(n639) );
  NAND2_X2 U473 ( .A1(n639), .A2(n516), .ZN(n272) );
  INV_X4 U474 ( .A(n272), .ZN(n709) );
  MUX2_X2 U475 ( .A(n512), .B(n91), .S(n709), .Z(n640) );
  INV_X4 U476 ( .A(n269), .ZN(n647) );
  NAND3_X2 U477 ( .A1(n195), .A2(n185), .A3(n252), .ZN(n665) );
  NOR3_X2 U478 ( .A1(n647), .A2(n641), .A3(n665), .ZN(n642) );
  MUX2_X2 U479 ( .A(n88), .B(n512), .S(n642), .Z(n643) );
  INV_X4 U480 ( .A(n644), .ZN(n646) );
  NAND2_X2 U481 ( .A1(n264), .A2(n191), .ZN(n181) );
  INV_X4 U482 ( .A(n181), .ZN(n648) );
  NAND3_X2 U483 ( .A1(n165), .A2(n649), .A3(n648), .ZN(n661) );
  INV_X4 U484 ( .A(n661), .ZN(n667) );
  NAND2_X2 U485 ( .A1(n650), .A2(n516), .ZN(n651) );
  NAND3_X2 U486 ( .A1(n651), .A2(n656), .A3(n706), .ZN(n314) );
  NAND4_X2 U487 ( .A1(n274), .A2(n329), .A3(n667), .A4(n676), .ZN(n327) );
  INV_X4 U488 ( .A(n327), .ZN(n652) );
  NAND2_X2 U489 ( .A1(n655), .A2(n652), .ZN(n653) );
  NAND2_X2 U490 ( .A1(n653), .A2(n516), .ZN(n328) );
  INV_X4 U491 ( .A(n328), .ZN(n715) );
  MUX2_X2 U492 ( .A(n512), .B(n84), .S(n715), .Z(n654) );
  INV_X4 U493 ( .A(n655), .ZN(n669) );
  NAND2_X2 U494 ( .A1(n669), .A2(n516), .ZN(n712) );
  INV_X4 U495 ( .A(n656), .ZN(n300) );
  NOR2_X2 U496 ( .A1(n300), .A2(n334), .ZN(n658) );
  INV_X4 U497 ( .A(n336), .ZN(n657) );
  NAND4_X2 U498 ( .A1(n658), .A2(n261), .A3(n657), .A4(n712), .ZN(n337) );
  INV_X4 U499 ( .A(n337), .ZN(n708) );
  MUX2_X2 U500 ( .A(n76), .B(n512), .S(n708), .Z(n660) );
  INV_X4 U501 ( .A(n329), .ZN(n719) );
  NOR3_X2 U502 ( .A1(n248), .A2(n719), .A3(n661), .ZN(n662) );
  NOR2_X2 U503 ( .A1(n517), .A2(n662), .ZN(n663) );
  MUX2_X2 U504 ( .A(n664), .B(WriteBus[120]), .S(n663), .Z(n483) );
  INV_X4 U505 ( .A(n665), .ZN(n668) );
  INV_X4 U506 ( .A(n334), .ZN(n666) );
  INV_X4 U507 ( .A(n706), .ZN(n286) );
  INV_X4 U508 ( .A(n193), .ZN(n696) );
  INV_X4 U509 ( .A(n265), .ZN(n698) );
  INV_X4 U510 ( .A(n284), .ZN(n699) );
  INV_X4 U511 ( .A(n232), .ZN(n700) );
  INV_X4 U512 ( .A(n169), .ZN(n701) );
  INV_X4 U513 ( .A(n268), .ZN(n702) );
  INV_X4 U514 ( .A(n220), .ZN(n704) );
  INV_X4 U515 ( .A(n330), .ZN(n707) );
  INV_X4 U516 ( .A(n270), .ZN(n710) );
  INV_X4 U517 ( .A(n333), .ZN(n711) );
  INV_X4 U518 ( .A(n313), .ZN(n713) );
  INV_X4 U519 ( .A(n353), .ZN(n714) );
  INV_X4 U520 ( .A(n326), .ZN(n716) );
  INV_X4 U521 ( .A(n206), .ZN(n717) );
  INV_X4 U522 ( .A(n163), .ZN(n718) );
endmodule


module Output_top ( clock, reset_n, start, CdfMin, divisor, M2SP_ReadBus, 
        M2SP_ReadAddress, M3SP_ReadBus, M3SP_ReadAddress, WriteEnable, 
        Output_MEMBus, Output_MEMAddress, done, output_base_offset );
  input [19:0] CdfMin;
  input [19:0] divisor;
  input [127:0] M2SP_ReadBus;
  output [15:0] M2SP_ReadAddress;
  input [127:0] M3SP_ReadBus;
  output [15:0] M3SP_ReadAddress;
  output [127:0] Output_MEMBus;
  output [15:0] Output_MEMAddress;
  input clock, reset_n, start, output_base_offset;
  output WriteEnable, done;
  wire   start_to_stage_two, start_to_stage_three, start_to_stage_four,
         start_to_stage_five, n15, n16;
  wire   [19:0] DataToStageThree;
  wire   [27:0] DataToStageFour;
  wire   [7:0] result;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  Output_Fetch_MEM stage1 ( .clock(clock), .reset_n(n15), .start(start), 
        .ReadBus(M3SP_ReadBus), .ReadAddress(M3SP_ReadAddress), .DataOut({
        M2SP_ReadAddress[15], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, M2SP_ReadAddress[7:0]}), .StartOut(
        start_to_stage_two), .output_base_offset(output_base_offset), .done(
        done) );
  Output_Fetch_Cdf stage2 ( .clock(clock), .reset_n(n15), .ReadBus(
        M2SP_ReadBus), .DataOut(DataToStageThree), .StartIn(start_to_stage_two), .StartOut(start_to_stage_three) );
  Output_TopExpression stage3 ( .clock(clock), .reset_n(n15), .DataIn(
        DataToStageThree), .CdfMin(CdfMin), .StartIn(start_to_stage_three), 
        .StartOut(start_to_stage_four), .DataOut(DataToStageFour) );
  Output_Result stage4 ( .clock(clock), .reset_n(n15), .DataIn(DataToStageFour), .StartIn(start_to_stage_four), .Divisor(divisor), .StartOut(
        start_to_stage_five), .DataOut(result) );
  Output_Store stage5 ( .clock(clock), .reset_n(n15), .StartIn(
        start_to_stage_five), .ResultIn(result), .WriteBus(Output_MEMBus), 
        .WriteAddress(Output_MEMAddress), .WriteEnable(WriteEnable), 
        .output_base_offset(output_base_offset) );
  INV_X4 U1 ( .A(1'b1), .ZN(M2SP_ReadAddress[8]) );
  INV_X4 U3 ( .A(1'b1), .ZN(M2SP_ReadAddress[9]) );
  INV_X4 U5 ( .A(1'b1), .ZN(M2SP_ReadAddress[10]) );
  INV_X4 U7 ( .A(1'b1), .ZN(M2SP_ReadAddress[11]) );
  INV_X4 U9 ( .A(1'b1), .ZN(M2SP_ReadAddress[12]) );
  INV_X4 U11 ( .A(1'b1), .ZN(M2SP_ReadAddress[13]) );
  INV_X4 U13 ( .A(1'b1), .ZN(M2SP_ReadAddress[14]) );
  INV_X4 U15 ( .A(n16), .ZN(n15) );
  INV_X4 U16 ( .A(reset_n), .ZN(n16) );
endmodule


module Controllor ( clock, reset_n, start, output_start, input_start, 
        input_done, output_done, Cdf_Min, Cdf_Min_Out, Divisor, 
        output_base_offset, input_base_offset, cdf_valid );
  input [19:0] Cdf_Min;
  output [19:0] Cdf_Min_Out;
  output [19:0] Divisor;
  input clock, reset_n, start, input_done, output_done, cdf_valid;
  output output_start, input_start, output_base_offset, input_base_offset;
  wire   \U3/U1/Z_0 , \U14/Z_1 , \U14/Z_2 , \U14/Z_3 , \U14/Z_4 , \U14/Z_5 ,
         \U14/Z_6 , \U14/Z_7 , \U14/Z_8 , \U14/Z_10 , \U14/Z_11 , \U14/Z_12 ,
         \U14/Z_13 , \U14/Z_14 , \U14/Z_15 , \U14/Z_16 , \U14/Z_17 ,
         \U14/Z_18 , \U14/Z_19 , \U13/DATA1_0 , \U11/DATA1_0 , \r311/DIFF[1] ,
         \r311/DIFF[2] , \r311/DIFF[3] , \r311/DIFF[4] , \r311/DIFF[5] ,
         \r311/DIFF[6] , \r311/DIFF[7] , \r311/DIFF[8] , \r311/DIFF[9] ,
         \r311/DIFF[10] , \r311/DIFF[11] , \r311/DIFF[12] , \r311/DIFF[13] ,
         \r311/DIFF[14] , \r311/DIFF[15] , \r311/DIFF[16] , \r311/DIFF[17] ,
         \r311/DIFF[18] , \r311/DIFF[19] , n27, n28, n29, n30, n31, n35, n36,
         n37, n42, n46, n47, n48, n51, n52, n54, n73, n75, n76, n79, n80, n81,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n280, n281, n282, n283,
         n284, n285, n286, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385;
  assign Cdf_Min_Out[0] = \U3/U1/Z_0 ;
  assign Cdf_Min_Out[1] = \U14/Z_1 ;
  assign Cdf_Min_Out[2] = \U14/Z_2 ;
  assign Cdf_Min_Out[3] = \U14/Z_3 ;
  assign Cdf_Min_Out[4] = \U14/Z_4 ;
  assign Cdf_Min_Out[5] = \U14/Z_5 ;
  assign Cdf_Min_Out[6] = \U14/Z_6 ;
  assign Cdf_Min_Out[7] = \U14/Z_7 ;
  assign Cdf_Min_Out[8] = \U14/Z_8 ;
  assign Cdf_Min_Out[10] = \U14/Z_10 ;
  assign Cdf_Min_Out[11] = \U14/Z_11 ;
  assign Cdf_Min_Out[12] = \U14/Z_12 ;
  assign Cdf_Min_Out[14] = \U14/Z_14 ;
  assign Cdf_Min_Out[15] = \U14/Z_15 ;
  assign Cdf_Min_Out[16] = \U14/Z_16 ;
  assign Cdf_Min_Out[17] = \U14/Z_17 ;
  assign Cdf_Min_Out[18] = \U14/Z_18 ;
  assign Cdf_Min_Out[19] = \U14/Z_19 ;
  assign \U13/DATA1_0  = input_done;
  assign \U11/DATA1_0  = start;
  assign Divisor[1] = \r311/DIFF[1] ;
  assign Divisor[2] = \r311/DIFF[2] ;
  assign Divisor[3] = \r311/DIFF[3] ;
  assign Divisor[4] = \r311/DIFF[4] ;
  assign Divisor[5] = \r311/DIFF[5] ;
  assign Divisor[6] = \r311/DIFF[6] ;
  assign Divisor[7] = \r311/DIFF[7] ;
  assign Divisor[8] = \r311/DIFF[8] ;
  assign Divisor[9] = \r311/DIFF[9] ;
  assign Divisor[10] = \r311/DIFF[10] ;
  assign Divisor[11] = \r311/DIFF[11] ;
  assign Divisor[12] = \r311/DIFF[12] ;
  assign Divisor[13] = \r311/DIFF[13] ;
  assign Divisor[14] = \r311/DIFF[14] ;
  assign Divisor[15] = \r311/DIFF[15] ;
  assign Divisor[16] = \r311/DIFF[16] ;
  assign Divisor[17] = \r311/DIFF[17] ;
  assign Divisor[18] = \r311/DIFF[18] ;
  assign Divisor[19] = \r311/DIFF[19] ;

  DFF_X2 RepeatState_reg ( .D(n131), .CK(clock), .QN(n126) );
  DFF_X1 \cdf_min1_reg[0]  ( .D(n123), .CK(cdf_valid), .Q(n177) );
  DFF_X1 \cdf_min1_reg[1]  ( .D(n122), .CK(cdf_valid), .Q(n192) );
  DFF_X1 \cdf_min1_reg[2]  ( .D(n121), .CK(cdf_valid), .Q(n206), .QN(n81) );
  DFF_X1 \cdf_min1_reg[3]  ( .D(n120), .CK(cdf_valid), .Q(n196), .QN(n80) );
  DFF_X1 \cdf_min1_reg[4]  ( .D(n119), .CK(cdf_valid), .Q(n195), .QN(n79) );
  DFF_X1 \cdf_min1_reg[5]  ( .D(n118), .CK(cdf_valid), .Q(n203) );
  DFF_X1 \cdf_min1_reg[6]  ( .D(n117), .CK(cdf_valid), .Q(n215) );
  DFF_X1 \cdf_min1_reg[7]  ( .D(n116), .CK(cdf_valid), .Q(n217), .QN(n76) );
  DFF_X1 \cdf_min1_reg[8]  ( .D(n115), .CK(cdf_valid), .Q(n193), .QN(n75) );
  DFF_X1 \cdf_min1_reg[9]  ( .D(n114), .CK(cdf_valid), .Q(n204) );
  DFF_X1 \cdf_min1_reg[10]  ( .D(n113), .CK(cdf_valid), .Q(n207), .QN(n73) );
  DFF_X1 \cdf_min1_reg[11]  ( .D(n112), .CK(cdf_valid), .Q(n205) );
  DFF_X1 \cdf_min1_reg[12]  ( .D(n111), .CK(n310), .Q(n210) );
  DFF_X1 \cdf_min1_reg[13]  ( .D(n110), .CK(cdf_valid), .Q(n211) );
  DFF_X1 \cdf_min1_reg[14]  ( .D(n109), .CK(n310), .Q(n212) );
  DFF_X1 \cdf_min1_reg[15]  ( .D(n108), .CK(n310), .Q(n213) );
  DFF_X1 \cdf_min1_reg[16]  ( .D(n107), .CK(cdf_valid), .Q(n214) );
  DFF_X1 \cdf_min1_reg[17]  ( .D(n106), .CK(n310), .Q(n209) );
  DFF_X1 \cdf_min1_reg[18]  ( .D(n105), .CK(cdf_valid), .Q(n187) );
  DFF_X1 \cdf_min1_reg[19]  ( .D(n104), .CK(n310), .Q(n188) );
  DFF_X1 \cdf_min0_reg[19]  ( .D(n103), .CK(cdf_valid), .Q(n179) );
  DFF_X1 \cdf_min0_reg[18]  ( .D(n102), .CK(n310), .Q(n178) );
  DFF_X1 \cdf_min0_reg[17]  ( .D(n101), .CK(cdf_valid), .Q(n186) );
  DFF_X1 \cdf_min0_reg[16]  ( .D(n100), .CK(n310), .Q(n201) );
  DFF_X1 \cdf_min0_reg[15]  ( .D(n99), .CK(cdf_valid), .Q(n200) );
  DFF_X1 \cdf_min0_reg[14]  ( .D(n98), .CK(n310), .Q(n199) );
  DFF_X1 \cdf_min0_reg[13]  ( .D(n97), .CK(cdf_valid), .Q(n198) );
  DFF_X1 \cdf_min0_reg[12]  ( .D(n96), .CK(n310), .Q(n208) );
  DFF_X1 \cdf_min0_reg[11]  ( .D(n95), .CK(n310), .Q(n185) );
  DFF_X1 \cdf_min0_reg[10]  ( .D(n94), .CK(n310), .Q(n194), .QN(n54) );
  DFF_X1 \cdf_min0_reg[9]  ( .D(n93), .CK(n310), .Q(n184) );
  DFF_X1 \cdf_min0_reg[8]  ( .D(n92), .CK(n310), .Q(n180), .QN(n52) );
  DFF_X1 \cdf_min0_reg[7]  ( .D(n91), .CK(n310), .Q(n216), .QN(n51) );
  DFF_X1 \cdf_min0_reg[6]  ( .D(n90), .CK(n310), .Q(n197) );
  DFF_X1 \cdf_min0_reg[5]  ( .D(n89), .CK(n310), .Q(n183) );
  DFF_X1 \cdf_min0_reg[4]  ( .D(n88), .CK(n310), .Q(n182), .QN(n48) );
  DFF_X1 \cdf_min0_reg[3]  ( .D(n87), .CK(n310), .Q(n190), .QN(n47) );
  DFF_X1 \cdf_min0_reg[2]  ( .D(n86), .CK(n310), .Q(n202), .QN(n46) );
  DFF_X1 \cdf_min0_reg[1]  ( .D(n85), .CK(n310), .Q(n181) );
  DFF_X1 \cdf_min0_reg[0]  ( .D(n84), .CK(n310), .Q(n191) );
  AND2_X1 U82 ( .A1(n30), .A2(n31), .ZN(n36) );
  OAI22_X2 U67 ( .A1(n189), .A2(n381), .B1(n27), .B2(n28), .ZN(n129) );
  OAI22_X2 U71 ( .A1(n31), .A2(n124), .B1(n29), .B2(n30), .ZN(n130) );
  NOR2_X2 U72 ( .A1(n382), .A2(n126), .ZN(n29) );
  OAI22_X2 U79 ( .A1(n42), .A2(n31), .B1(n37), .B2(n384), .ZN(n132) );
  NAND2_X2 U83 ( .A1(n127), .A2(n384), .ZN(n31) );
  NAND2_X2 U84 ( .A1(n384), .A2(n383), .ZN(n30) );
  DFFR_X2 output_base_offset_reg ( .D(n128), .CK(clock), .RN(n314), .Q(n237), 
        .QN(n306) );
  DFFR_X2 output_start_reg ( .D(n130), .CK(clock), .RN(n314), .Q(output_start), 
        .QN(n124) );
  DFFR_X2 input_start_reg ( .D(n132), .CK(clock), .RN(n314), .Q(input_start), 
        .QN(n42) );
  DFFR_X2 input_base_offset_reg ( .D(n129), .CK(clock), .RN(n314), .Q(
        input_base_offset), .QN(n189) );
  DFFR_X2 \State_reg[0]  ( .D(n134), .CK(clock), .RN(reset_n), .Q(n383), .QN(
        n127) );
  DFFR_X2 \State_reg[1]  ( .D(n133), .CK(clock), .RN(n314), .Q(n384) );
  NAND2_X1 U3 ( .A1(n375), .A2(n374), .ZN(n285) );
  NAND2_X2 U4 ( .A1(n293), .A2(n294), .ZN(\U14/Z_15 ) );
  INV_X4 U5 ( .A(n319), .ZN(\U14/Z_1 ) );
  NOR2_X2 U6 ( .A1(n370), .A2(\U14/Z_16 ), .ZN(n371) );
  NOR2_X2 U7 ( .A1(output_base_offset), .A2(n180), .ZN(n256) );
  NAND2_X2 U8 ( .A1(n297), .A2(n298), .ZN(\U14/Z_12 ) );
  INV_X4 U9 ( .A(n312), .ZN(n282) );
  INV_X8 U10 ( .A(n282), .ZN(output_base_offset) );
  NOR2_X2 U11 ( .A1(\U14/Z_14 ), .A2(n174), .ZN(n225) );
  NAND2_X1 U12 ( .A1(n271), .A2(n305), .ZN(n174) );
  INV_X2 U13 ( .A(n320), .ZN(n351) );
  NAND3_X2 U14 ( .A1(n328), .A2(n348), .A3(n337), .ZN(n175) );
  NAND3_X1 U15 ( .A1(n333), .A2(n276), .A3(n331), .ZN(n176) );
  OR2_X1 U16 ( .A1(n206), .A2(n313), .ZN(n281) );
  INV_X4 U17 ( .A(n349), .ZN(\U14/Z_4 ) );
  INV_X1 U18 ( .A(n337), .ZN(n338) );
  INV_X4 U19 ( .A(\U14/Z_15 ), .ZN(n247) );
  INV_X2 U20 ( .A(n340), .ZN(n341) );
  INV_X1 U21 ( .A(n359), .ZN(n363) );
  NAND2_X2 U22 ( .A1(n327), .A2(n219), .ZN(n220) );
  NAND2_X2 U23 ( .A1(n218), .A2(\U14/Z_6 ), .ZN(n221) );
  NAND2_X2 U24 ( .A1(n220), .A2(n221), .ZN(\r311/DIFF[6] ) );
  INV_X4 U25 ( .A(n327), .ZN(n218) );
  INV_X4 U26 ( .A(\U14/Z_6 ), .ZN(n219) );
  INV_X1 U27 ( .A(n348), .ZN(\U14/Z_6 ) );
  NAND2_X2 U28 ( .A1(n194), .A2(n292), .ZN(n222) );
  NAND2_X1 U29 ( .A1(n207), .A2(n312), .ZN(n223) );
  NAND2_X2 U30 ( .A1(n222), .A2(n223), .ZN(\U14/Z_10 ) );
  NAND2_X1 U31 ( .A1(\U14/Z_10 ), .A2(n335), .ZN(n243) );
  XNOR2_X2 U32 ( .A(n224), .B(\U14/Z_2 ), .ZN(\r311/DIFF[2] ) );
  AND2_X4 U33 ( .A1(n317), .A2(n319), .ZN(n224) );
  NOR2_X2 U34 ( .A1(n225), .A2(n362), .ZN(n245) );
  OAI22_X1 U35 ( .A1(n360), .A2(n361), .B1(n305), .B2(n373), .ZN(n362) );
  NAND2_X1 U36 ( .A1(n176), .A2(n336), .ZN(n269) );
  INV_X4 U37 ( .A(n231), .ZN(n232) );
  INV_X2 U38 ( .A(n357), .ZN(n356) );
  INV_X1 U39 ( .A(n318), .ZN(\U14/Z_2 ) );
  INV_X2 U40 ( .A(n344), .ZN(\U14/Z_3 ) );
  INV_X4 U41 ( .A(n320), .ZN(n226) );
  NOR2_X2 U42 ( .A1(n312), .A2(n197), .ZN(n229) );
  NAND2_X2 U43 ( .A1(\U14/Z_17 ), .A2(n376), .ZN(n286) );
  XNOR2_X2 U44 ( .A(n226), .B(\U14/Z_3 ), .ZN(\r311/DIFF[3] ) );
  INV_X2 U45 ( .A(n228), .ZN(n348) );
  INV_X4 U46 ( .A(n326), .ZN(n328) );
  NOR2_X2 U47 ( .A1(n229), .A2(n230), .ZN(n228) );
  OR2_X2 U48 ( .A1(n377), .A2(\U14/Z_18 ), .ZN(n263) );
  NAND2_X2 U49 ( .A1(n377), .A2(\U14/Z_18 ), .ZN(n262) );
  INV_X4 U50 ( .A(n364), .ZN(n369) );
  INV_X1 U51 ( .A(n337), .ZN(\U14/Z_5 ) );
  INV_X4 U52 ( .A(n321), .ZN(n252) );
  NAND2_X1 U53 ( .A1(n378), .A2(\U14/Z_19 ), .ZN(n274) );
  NAND2_X2 U54 ( .A1(n198), .A2(n282), .ZN(n299) );
  INV_X4 U55 ( .A(n368), .ZN(n305) );
  NAND2_X1 U56 ( .A1(n305), .A2(n373), .ZN(n360) );
  INV_X1 U57 ( .A(n336), .ZN(Cdf_Min_Out[9]) );
  NOR2_X1 U58 ( .A1(n215), .A2(n313), .ZN(n230) );
  AOI21_X4 U59 ( .B1(n347), .B2(n346), .A(n345), .ZN(n352) );
  XOR2_X2 U60 ( .A(n271), .B(\U14/Z_11 ), .Z(\r311/DIFF[11] ) );
  NAND2_X1 U61 ( .A1(n373), .A2(n372), .ZN(n231) );
  NAND2_X2 U62 ( .A1(n232), .A2(n365), .ZN(n366) );
  NAND2_X2 U63 ( .A1(n359), .A2(\U14/Z_12 ), .ZN(n233) );
  NAND2_X1 U64 ( .A1(n359), .A2(\U14/Z_12 ), .ZN(n234) );
  NAND2_X2 U65 ( .A1(n359), .A2(\U14/Z_12 ), .ZN(n357) );
  NOR2_X2 U66 ( .A1(n308), .A2(n247), .ZN(n235) );
  NOR2_X2 U68 ( .A1(n369), .A2(n236), .ZN(n370) );
  INV_X4 U69 ( .A(n235), .ZN(n236) );
  NAND2_X2 U70 ( .A1(n226), .A2(n344), .ZN(n321) );
  NAND2_X2 U73 ( .A1(n376), .A2(n375), .ZN(n377) );
  NOR2_X4 U74 ( .A1(n312), .A2(n190), .ZN(n290) );
  INV_X4 U75 ( .A(n175), .ZN(n333) );
  INV_X1 U76 ( .A(\U14/Z_12 ), .ZN(n354) );
  NAND2_X1 U77 ( .A1(\U14/Z_12 ), .A2(\U14/Z_13 ), .ZN(n308) );
  NAND2_X1 U78 ( .A1(n234), .A2(n355), .ZN(\r311/DIFF[12] ) );
  XOR2_X2 U80 ( .A(n329), .B(\U14/Z_7 ), .Z(\r311/DIFF[7] ) );
  NAND2_X2 U81 ( .A1(n271), .A2(n305), .ZN(n365) );
  OR2_X4 U85 ( .A1(n312), .A2(n202), .ZN(n280) );
  NOR2_X2 U86 ( .A1(n312), .A2(n325), .ZN(n277) );
  NAND2_X1 U87 ( .A1(n208), .A2(n313), .ZN(n297) );
  INV_X2 U88 ( .A(n342), .ZN(n343) );
  NOR2_X1 U89 ( .A1(n313), .A2(n324), .ZN(n278) );
  INV_X2 U90 ( .A(n237), .ZN(n238) );
  INV_X4 U91 ( .A(n317), .ZN(\U3/U1/Z_0 ) );
  INV_X2 U92 ( .A(n366), .ZN(n246) );
  NAND2_X2 U93 ( .A1(n201), .A2(n282), .ZN(n239) );
  NAND2_X1 U94 ( .A1(n214), .A2(n312), .ZN(n240) );
  NAND2_X2 U95 ( .A1(n239), .A2(n240), .ZN(\U14/Z_16 ) );
  NOR2_X2 U96 ( .A1(Cdf_Min_Out[13]), .A2(n356), .ZN(n289) );
  NOR2_X2 U97 ( .A1(\U14/Z_4 ), .A2(n228), .ZN(n350) );
  NAND2_X2 U98 ( .A1(n312), .A2(n76), .ZN(n342) );
  NOR2_X2 U99 ( .A1(n313), .A2(n196), .ZN(n291) );
  NAND2_X2 U100 ( .A1(n369), .A2(n361), .ZN(n359) );
  NAND2_X2 U101 ( .A1(n242), .A2(n241), .ZN(n244) );
  NAND2_X2 U102 ( .A1(n244), .A2(n243), .ZN(\r311/DIFF[10] ) );
  INV_X2 U103 ( .A(\U14/Z_10 ), .ZN(n241) );
  INV_X2 U104 ( .A(n335), .ZN(n242) );
  NOR2_X2 U105 ( .A1(Cdf_Min_Out[9]), .A2(n176), .ZN(n335) );
  NAND2_X2 U106 ( .A1(n245), .A2(n267), .ZN(\r311/DIFF[14] ) );
  NAND2_X2 U107 ( .A1(n246), .A2(n247), .ZN(n248) );
  NAND2_X2 U108 ( .A1(n248), .A2(n367), .ZN(\r311/DIFF[15] ) );
  NAND2_X2 U109 ( .A1(n330), .A2(n332), .ZN(n250) );
  NAND2_X2 U110 ( .A1(n249), .A2(\U14/Z_8 ), .ZN(n251) );
  NAND2_X2 U111 ( .A1(n250), .A2(n251), .ZN(\r311/DIFF[8] ) );
  INV_X4 U112 ( .A(n330), .ZN(n249) );
  NAND2_X2 U113 ( .A1(n321), .A2(n253), .ZN(n254) );
  NAND2_X2 U114 ( .A1(n252), .A2(\U14/Z_4 ), .ZN(n255) );
  NAND2_X2 U115 ( .A1(n254), .A2(n255), .ZN(\r311/DIFF[4] ) );
  INV_X1 U116 ( .A(\U14/Z_4 ), .ZN(n253) );
  NOR2_X1 U117 ( .A1(n193), .A2(n292), .ZN(n257) );
  OR2_X4 U118 ( .A1(n256), .A2(n257), .ZN(n332) );
  NAND2_X1 U119 ( .A1(n326), .A2(n259), .ZN(n260) );
  NAND2_X2 U120 ( .A1(n258), .A2(\U14/Z_5 ), .ZN(n261) );
  NAND2_X2 U121 ( .A1(n260), .A2(n261), .ZN(\r311/DIFF[5] ) );
  INV_X1 U122 ( .A(n326), .ZN(n258) );
  INV_X1 U123 ( .A(\U14/Z_5 ), .ZN(n259) );
  NAND2_X2 U124 ( .A1(n263), .A2(n262), .ZN(\r311/DIFF[18] ) );
  NAND2_X1 U125 ( .A1(\U14/Z_1 ), .A2(n264), .ZN(n265) );
  NAND2_X1 U126 ( .A1(n319), .A2(\U3/U1/Z_0 ), .ZN(n266) );
  NAND2_X2 U127 ( .A1(n265), .A2(n266), .ZN(\r311/DIFF[1] ) );
  INV_X1 U128 ( .A(\U3/U1/Z_0 ), .ZN(n264) );
  NAND2_X1 U129 ( .A1(n363), .A2(\U14/Z_14 ), .ZN(n267) );
  NAND2_X2 U130 ( .A1(n283), .A2(n284), .ZN(\U14/Z_14 ) );
  NAND2_X2 U131 ( .A1(n268), .A2(n339), .ZN(n270) );
  NAND2_X2 U132 ( .A1(n269), .A2(n270), .ZN(\r311/DIFF[9] ) );
  INV_X4 U133 ( .A(n334), .ZN(n268) );
  NAND2_X1 U134 ( .A1(n333), .A2(n331), .ZN(n330) );
  INV_X4 U135 ( .A(n344), .ZN(n345) );
  OAI22_X2 U136 ( .A1(n312), .A2(n184), .B1(n238), .B2(n204), .ZN(n336) );
  INV_X4 U137 ( .A(n336), .ZN(n339) );
  XNOR2_X2 U138 ( .A(n367), .B(\U14/Z_16 ), .ZN(\r311/DIFF[16] ) );
  INV_X16 U139 ( .A(n313), .ZN(n312) );
  OR2_X2 U140 ( .A1(n277), .A2(n278), .ZN(n326) );
  OAI22_X2 U141 ( .A1(n312), .A2(n182), .B1(n195), .B2(n313), .ZN(n349) );
  INV_X16 U142 ( .A(n307), .ZN(n313) );
  NAND3_X2 U143 ( .A1(n302), .A2(n352), .A3(n351), .ZN(n271) );
  NAND2_X2 U144 ( .A1(n272), .A2(n273), .ZN(n275) );
  NAND2_X2 U145 ( .A1(n275), .A2(n274), .ZN(\r311/DIFF[19] ) );
  INV_X2 U146 ( .A(n378), .ZN(n272) );
  INV_X2 U147 ( .A(\U14/Z_19 ), .ZN(n273) );
  OAI22_X2 U148 ( .A1(output_base_offset), .A2(n180), .B1(n193), .B2(n282), 
        .ZN(n276) );
  NAND2_X2 U149 ( .A1(n280), .A2(n281), .ZN(n318) );
  OAI22_X2 U150 ( .A1(n312), .A2(n191), .B1(n313), .B2(n177), .ZN(n317) );
  OAI22_X2 U151 ( .A1(n312), .A2(n183), .B1(n313), .B2(n203), .ZN(n337) );
  OAI22_X2 U152 ( .A1(n312), .A2(n181), .B1(n313), .B2(n192), .ZN(n319) );
  NAND2_X2 U153 ( .A1(n199), .A2(n282), .ZN(n283) );
  NAND2_X1 U154 ( .A1(n212), .A2(output_base_offset), .ZN(n284) );
  NAND2_X2 U155 ( .A1(n285), .A2(n286), .ZN(\r311/DIFF[17] ) );
  INV_X4 U156 ( .A(n358), .ZN(Cdf_Min_Out[13]) );
  INV_X1 U157 ( .A(\U14/Z_13 ), .ZN(n358) );
  OR2_X1 U158 ( .A1(n247), .A2(n373), .ZN(n295) );
  NOR2_X2 U159 ( .A1(n358), .A2(n233), .ZN(n288) );
  OR2_X2 U160 ( .A1(n288), .A2(n289), .ZN(\r311/DIFF[13] ) );
  OR2_X2 U161 ( .A1(n290), .A2(n291), .ZN(n344) );
  NAND2_X2 U162 ( .A1(n200), .A2(n292), .ZN(n293) );
  NAND2_X1 U163 ( .A1(n213), .A2(n312), .ZN(n294) );
  INV_X1 U164 ( .A(n312), .ZN(n292) );
  OR2_X1 U165 ( .A1(n247), .A2(n372), .ZN(n296) );
  NAND3_X2 U166 ( .A1(n371), .A2(n296), .A3(n295), .ZN(n374) );
  NAND2_X1 U167 ( .A1(n210), .A2(n312), .ZN(n298) );
  NAND2_X1 U168 ( .A1(n211), .A2(n312), .ZN(n300) );
  NAND2_X2 U169 ( .A1(n299), .A2(n300), .ZN(\U14/Z_13 ) );
  NAND2_X2 U170 ( .A1(n353), .A2(n350), .ZN(n301) );
  NAND3_X2 U171 ( .A1(n302), .A2(n352), .A3(n351), .ZN(n364) );
  INV_X4 U172 ( .A(n301), .ZN(n302) );
  INV_X4 U173 ( .A(input_base_offset), .ZN(n309) );
  OAI21_X2 U174 ( .B1(n29), .B2(n30), .A(n31), .ZN(n27) );
  INV_X4 U175 ( .A(n315), .ZN(n314) );
  INV_X4 U176 ( .A(reset_n), .ZN(n315) );
  INV_X4 U177 ( .A(n311), .ZN(n310) );
  INV_X4 U178 ( .A(cdf_valid), .ZN(n311) );
  AOI22_X2 U179 ( .A1(\U11/DATA1_0 ), .A2(n127), .B1(n380), .B2(n383), .ZN(n37) );
  OAI21_X2 U180 ( .B1(n385), .B2(n384), .A(n127), .ZN(n134) );
  OAI21_X2 U181 ( .B1(n127), .B2(n380), .A(n36), .ZN(n133) );
  OR2_X1 U182 ( .A1(n35), .A2(n303), .ZN(n131) );
  AND3_X4 U183 ( .A1(\U13/DATA1_0 ), .A2(n379), .A3(n314), .ZN(n303) );
  AOI21_X2 U184 ( .B1(n314), .B2(n36), .A(n126), .ZN(n35) );
  INV_X1 U185 ( .A(n264), .ZN(Divisor[0]) );
  NAND2_X2 U186 ( .A1(\U14/Z_11 ), .A2(n305), .ZN(n372) );
  NAND2_X1 U187 ( .A1(n51), .A2(n238), .ZN(n340) );
  NOR2_X1 U188 ( .A1(output_base_offset), .A2(n30), .ZN(n316) );
  NAND2_X1 U189 ( .A1(n328), .A2(n337), .ZN(n327) );
  NAND3_X1 U190 ( .A1(n369), .A2(n354), .A3(n361), .ZN(n355) );
  NAND2_X2 U191 ( .A1(\U14/Z_12 ), .A2(\U14/Z_13 ), .ZN(n368) );
  INV_X4 U192 ( .A(n306), .ZN(n307) );
  INV_X4 U193 ( .A(n30), .ZN(n379) );
  INV_X4 U194 ( .A(n27), .ZN(n381) );
  NAND2_X2 U195 ( .A1(n189), .A2(n379), .ZN(n28) );
  MUX2_X2 U196 ( .A(output_base_offset), .B(n316), .S(n381), .Z(n128) );
  MUX2_X2 U197 ( .A(Cdf_Min[0]), .B(n177), .S(n189), .Z(n123) );
  MUX2_X2 U198 ( .A(n191), .B(Cdf_Min[0]), .S(n309), .Z(n84) );
  MUX2_X2 U199 ( .A(Cdf_Min[1]), .B(n192), .S(n309), .Z(n122) );
  MUX2_X2 U200 ( .A(n181), .B(Cdf_Min[1]), .S(n309), .Z(n85) );
  MUX2_X2 U201 ( .A(Cdf_Min[2]), .B(n206), .S(n309), .Z(n121) );
  MUX2_X2 U202 ( .A(n202), .B(Cdf_Min[2]), .S(n309), .Z(n86) );
  MUX2_X2 U203 ( .A(Cdf_Min[3]), .B(n196), .S(n309), .Z(n120) );
  MUX2_X2 U204 ( .A(n190), .B(Cdf_Min[3]), .S(n309), .Z(n87) );
  NAND3_X2 U205 ( .A1(n318), .A2(n319), .A3(n317), .ZN(n320) );
  MUX2_X2 U206 ( .A(Cdf_Min[4]), .B(n195), .S(n309), .Z(n119) );
  MUX2_X2 U207 ( .A(n182), .B(Cdf_Min[4]), .S(n309), .Z(n88) );
  MUX2_X2 U208 ( .A(Cdf_Min[5]), .B(n203), .S(n309), .Z(n118) );
  MUX2_X2 U209 ( .A(n183), .B(Cdf_Min[5]), .S(n309), .Z(n89) );
  NAND3_X2 U210 ( .A1(n46), .A2(n48), .A3(n47), .ZN(n322) );
  NOR3_X2 U211 ( .A1(n322), .A2(n181), .A3(n191), .ZN(n325) );
  NAND3_X2 U212 ( .A1(n81), .A2(n79), .A3(n80), .ZN(n323) );
  NOR3_X2 U213 ( .A1(n323), .A2(n192), .A3(n177), .ZN(n324) );
  MUX2_X2 U214 ( .A(Cdf_Min[6]), .B(n215), .S(n309), .Z(n117) );
  MUX2_X2 U215 ( .A(n197), .B(Cdf_Min[6]), .S(n309), .Z(n90) );
  MUX2_X2 U216 ( .A(Cdf_Min[7]), .B(n217), .S(n309), .Z(n116) );
  MUX2_X2 U217 ( .A(n216), .B(Cdf_Min[7]), .S(n309), .Z(n91) );
  NAND3_X2 U218 ( .A1(n328), .A2(n348), .A3(n337), .ZN(n329) );
  NAND2_X2 U219 ( .A1(n340), .A2(n342), .ZN(n331) );
  INV_X4 U220 ( .A(n331), .ZN(\U14/Z_7 ) );
  MUX2_X2 U221 ( .A(Cdf_Min[8]), .B(n193), .S(n309), .Z(n115) );
  MUX2_X2 U222 ( .A(n180), .B(Cdf_Min[8]), .S(n309), .Z(n92) );
  INV_X4 U223 ( .A(n332), .ZN(\U14/Z_8 ) );
  MUX2_X2 U224 ( .A(Cdf_Min[9]), .B(n204), .S(n309), .Z(n114) );
  MUX2_X2 U225 ( .A(n184), .B(Cdf_Min[9]), .S(n309), .Z(n93) );
  NAND3_X2 U226 ( .A1(n333), .A2(n276), .A3(n331), .ZN(n334) );
  MUX2_X2 U227 ( .A(n194), .B(Cdf_Min[10]), .S(n309), .Z(n94) );
  MUX2_X2 U228 ( .A(Cdf_Min[10]), .B(n207), .S(n309), .Z(n113) );
  MUX2_X2 U229 ( .A(Cdf_Min[11]), .B(n205), .S(n309), .Z(n112) );
  MUX2_X2 U230 ( .A(n185), .B(Cdf_Min[11]), .S(n309), .Z(n95) );
  NOR2_X2 U231 ( .A1(n338), .A2(n339), .ZN(n353) );
  NAND3_X2 U232 ( .A1(n54), .A2(n341), .A3(n52), .ZN(n347) );
  NAND3_X2 U233 ( .A1(n73), .A2(n343), .A3(n75), .ZN(n346) );
  OAI22_X2 U234 ( .A1(output_base_offset), .A2(n185), .B1(n205), .B2(n282), 
        .ZN(n361) );
  INV_X4 U235 ( .A(n361), .ZN(\U14/Z_11 ) );
  MUX2_X2 U236 ( .A(n208), .B(Cdf_Min[12]), .S(n309), .Z(n96) );
  MUX2_X2 U237 ( .A(Cdf_Min[12]), .B(n210), .S(n309), .Z(n111) );
  MUX2_X2 U238 ( .A(n198), .B(Cdf_Min[13]), .S(n309), .Z(n97) );
  MUX2_X2 U239 ( .A(Cdf_Min[13]), .B(n211), .S(n309), .Z(n110) );
  MUX2_X2 U240 ( .A(n199), .B(Cdf_Min[14]), .S(n309), .Z(n98) );
  MUX2_X2 U241 ( .A(Cdf_Min[14]), .B(n212), .S(n309), .Z(n109) );
  INV_X4 U242 ( .A(\U14/Z_14 ), .ZN(n373) );
  MUX2_X2 U243 ( .A(n200), .B(Cdf_Min[15]), .S(n309), .Z(n99) );
  MUX2_X2 U244 ( .A(Cdf_Min[15]), .B(n213), .S(n309), .Z(n108) );
  NAND2_X2 U245 ( .A1(n366), .A2(\U14/Z_15 ), .ZN(n367) );
  MUX2_X2 U246 ( .A(n201), .B(Cdf_Min[16]), .S(n309), .Z(n100) );
  MUX2_X2 U247 ( .A(Cdf_Min[16]), .B(n214), .S(n309), .Z(n107) );
  MUX2_X2 U248 ( .A(n186), .B(Cdf_Min[17]), .S(n309), .Z(n101) );
  MUX2_X2 U249 ( .A(Cdf_Min[17]), .B(n209), .S(n309), .Z(n106) );
  MUX2_X2 U250 ( .A(n186), .B(n209), .S(output_base_offset), .Z(\U14/Z_17 ) );
  INV_X4 U251 ( .A(\U14/Z_17 ), .ZN(n375) );
  INV_X4 U252 ( .A(n374), .ZN(n376) );
  MUX2_X2 U253 ( .A(n178), .B(Cdf_Min[18]), .S(n309), .Z(n102) );
  MUX2_X2 U254 ( .A(Cdf_Min[18]), .B(n187), .S(n309), .Z(n105) );
  MUX2_X2 U255 ( .A(n178), .B(n187), .S(output_base_offset), .Z(\U14/Z_18 ) );
  MUX2_X2 U256 ( .A(n179), .B(Cdf_Min[19]), .S(n309), .Z(n103) );
  MUX2_X2 U257 ( .A(Cdf_Min[19]), .B(n188), .S(n309), .Z(n104) );
  NAND2_X2 U258 ( .A1(\U14/Z_18 ), .A2(n377), .ZN(n378) );
  MUX2_X2 U259 ( .A(n179), .B(n188), .S(output_base_offset), .Z(\U14/Z_19 ) );
  INV_X4 U260 ( .A(\U13/DATA1_0 ), .ZN(n380) );
  INV_X4 U261 ( .A(output_done), .ZN(n382) );
  INV_X4 U262 ( .A(\U11/DATA1_0 ), .ZN(n385) );
endmodule


module Cdf_Fetch ( clock, reset_n, start, ReadBus, ReadAddr, AccumlateOut, 
        StartOut, StoreAddress, input_base_offset, done );
  input [127:0] ReadBus;
  output [15:0] ReadAddr;
  output [19:0] AccumlateOut;
  output [15:0] StoreAddress;
  input clock, reset_n, start, input_base_offset;
  output StartOut, done;
  wire   n208, n210, \U3/U1/DATA1_1 , \U3/U1/DATA1_2 , \U3/U1/DATA1_3 ,
         \U3/U1/DATA1_4 , \U3/U1/DATA1_5 , \U3/U1/DATA1_6 , \U3/U1/DATA1_7 ,
         \U8/DATA1_0 , \U8/DATA1_1 , \U8/DATA1_2 , \U8/DATA1_3 , \U8/DATA1_4 ,
         \U8/DATA1_5 , \U8/DATA1_6 , \U8/DATA1_7 , \U8/DATA1_8 , \U8/DATA1_9 ,
         \U8/DATA1_10 , \U8/DATA1_11 , \U8/DATA1_12 , \U8/DATA1_13 ,
         \U8/DATA1_14 , \U8/DATA1_15 , \U8/DATA1_16 , \U8/DATA1_17 ,
         \U8/DATA1_18 , \U8/DATA1_19 , \U7/Z_0 , \U7/Z_1 , \U7/Z_2 , \U7/Z_3 ,
         \U7/Z_4 , \U7/Z_5 , \U7/Z_6 , \U7/Z_7 , \U7/Z_8 , \U7/Z_9 , \U7/Z_10 ,
         \U7/Z_11 , \U7/Z_12 , \U7/Z_13 , \U7/Z_14 , \U7/Z_15 , \U7/Z_16 ,
         \U7/Z_17 , \U7/Z_18 , \U7/Z_19 , \U5/Z_0 , \U5/Z_1 , \U5/Z_2 ,
         \U5/Z_3 , \U5/Z_4 , \U5/Z_5 , \U5/Z_6 , \U5/Z_7 , \U5/Z_8 , \U5/Z_9 ,
         \U5/Z_10 , \U5/Z_11 , \U5/Z_12 , \U5/Z_13 , \U5/Z_14 , \U4/Z_0 ,
         \U4/DATA3_0 , \add_63/carry[8] , \add_63/carry[7] , \add_63/carry[6] ,
         \add_63/carry[5] , \add_63/carry[4] , \add_63/carry[3] ,
         \add_63/carry[2] , \add_63/A[0] , \add_63/A[1] , \add_63/A[2] ,
         \add_63/A[3] , \add_63/A[4] , \add_63/A[5] , \add_63/A[6] ,
         \add_63/A[7] , \add_63/A[8] , \add_60/A[0] , \add_60/A[1] ,
         \add_60/A[2] , \add_60/A[3] , \add_60/A[4] , \add_60/A[5] ,
         \add_60/A[6] , \add_60/A[7] , \add_60/A[8] , \add_60/A[9] ,
         \add_60/A[10] , \add_60/A[11] , \add_60/A[12] , \add_60/A[13] ,
         \add_60/A[14] , \add_60/A[15] , n1, n2, n4, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n26, n27, n28, n29, n30, n31, n32, n33, n34, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440;
  assign \U8/DATA1_0  = ReadBus[0];
  assign \U8/DATA1_1  = ReadBus[1];
  assign \U8/DATA1_2  = ReadBus[2];
  assign \U8/DATA1_3  = ReadBus[3];
  assign \U8/DATA1_4  = ReadBus[4];
  assign \U8/DATA1_5  = ReadBus[5];
  assign \U8/DATA1_6  = ReadBus[6];
  assign \U8/DATA1_7  = ReadBus[7];
  assign \U8/DATA1_8  = ReadBus[8];
  assign \U8/DATA1_9  = ReadBus[9];
  assign \U8/DATA1_10  = ReadBus[10];
  assign \U8/DATA1_11  = ReadBus[11];
  assign \U8/DATA1_12  = ReadBus[12];
  assign \U8/DATA1_13  = ReadBus[13];
  assign \U8/DATA1_14  = ReadBus[14];
  assign \U8/DATA1_15  = ReadBus[15];
  assign \U8/DATA1_16  = ReadBus[16];
  assign \U8/DATA1_17  = ReadBus[17];
  assign \U8/DATA1_18  = ReadBus[18];
  assign \U8/DATA1_19  = ReadBus[19];
  assign \U4/DATA3_0  = input_base_offset;

  HA_X1 \add_63/U1_1_1  ( .A(\add_63/A[1] ), .B(\add_63/A[0] ), .CO(
        \add_63/carry[2] ), .S(\U3/U1/DATA1_1 ) );
  HA_X1 \add_63/U1_1_2  ( .A(\add_63/A[2] ), .B(\add_63/carry[2] ), .CO(
        \add_63/carry[3] ), .S(\U3/U1/DATA1_2 ) );
  HA_X1 \add_63/U1_1_3  ( .A(\add_63/A[3] ), .B(\add_63/carry[3] ), .CO(
        \add_63/carry[4] ), .S(\U3/U1/DATA1_3 ) );
  HA_X1 \add_63/U1_1_4  ( .A(\add_63/A[4] ), .B(\add_63/carry[4] ), .CO(
        \add_63/carry[5] ), .S(\U3/U1/DATA1_4 ) );
  HA_X1 \add_63/U1_1_5  ( .A(\add_63/A[5] ), .B(\add_63/carry[5] ), .CO(
        \add_63/carry[6] ), .S(\U3/U1/DATA1_5 ) );
  HA_X1 \add_63/U1_1_6  ( .A(\add_63/A[6] ), .B(\add_63/carry[6] ), .CO(
        \add_63/carry[7] ), .S(\U3/U1/DATA1_6 ) );
  HA_X1 \add_63/U1_1_7  ( .A(\add_63/A[7] ), .B(\add_63/carry[7] ), .CO(
        \add_63/carry[8] ), .S(\U3/U1/DATA1_7 ) );
  SDFFR_X2 StartOut_reg ( .D(1'b0), .SI(start), .SE(n1), .CK(clock), .RN(
        reset_n), .Q(StartOut) );
  SDFFR_X2 done0_reg ( .D(1'b0), .SI(start), .SE(\add_63/A[8] ), .CK(clock), 
        .RN(reset_n), .Q(n210) );
  TBUF_X2 \ReadAddr_tri[0]  ( .A(\add_60/A[0] ), .EN(n395), .Z(ReadAddr[0]) );
  TBUF_X2 \ReadAddr_tri[1]  ( .A(\add_60/A[1] ), .EN(n395), .Z(ReadAddr[1]) );
  TBUF_X2 \ReadAddr_tri[2]  ( .A(\add_60/A[2] ), .EN(n395), .Z(ReadAddr[2]) );
  TBUF_X2 \ReadAddr_tri[3]  ( .A(\add_60/A[3] ), .EN(n395), .Z(ReadAddr[3]) );
  TBUF_X2 \ReadAddr_tri[4]  ( .A(\add_60/A[4] ), .EN(n395), .Z(ReadAddr[4]) );
  TBUF_X2 \ReadAddr_tri[5]  ( .A(\add_60/A[5] ), .EN(n395), .Z(ReadAddr[5]) );
  TBUF_X2 \ReadAddr_tri[6]  ( .A(\add_60/A[6] ), .EN(n395), .Z(ReadAddr[6]) );
  TBUF_X2 \ReadAddr_tri[7]  ( .A(\add_60/A[7] ), .EN(n395), .Z(ReadAddr[7]) );
  TBUF_X2 \ReadAddr_tri[8]  ( .A(\add_60/A[8] ), .EN(n395), .Z(ReadAddr[8]) );
  TBUF_X2 \ReadAddr_tri[9]  ( .A(\add_60/A[9] ), .EN(n395), .Z(ReadAddr[9]) );
  TBUF_X2 \ReadAddr_tri[10]  ( .A(\add_60/A[10] ), .EN(n395), .Z(ReadAddr[10])
         );
  TBUF_X2 \ReadAddr_tri[11]  ( .A(\add_60/A[11] ), .EN(n395), .Z(ReadAddr[11])
         );
  TBUF_X2 \ReadAddr_tri[12]  ( .A(\add_60/A[12] ), .EN(n395), .Z(ReadAddr[12])
         );
  TBUF_X2 \ReadAddr_tri[13]  ( .A(\add_60/A[13] ), .EN(n395), .Z(ReadAddr[13])
         );
  TBUF_X2 \ReadAddr_tri[14]  ( .A(\add_60/A[14] ), .EN(n395), .Z(ReadAddr[14])
         );
  TBUF_X2 \ReadAddr_tri[15]  ( .A(\add_60/A[15] ), .EN(n395), .Z(ReadAddr[15])
         );
  AND2_X1 U30 ( .A1(\U8/DATA1_19 ), .A2(n374), .ZN(\U7/Z_19 ) );
  AND2_X1 U31 ( .A1(\U8/DATA1_18 ), .A2(n374), .ZN(\U7/Z_18 ) );
  AND2_X1 U32 ( .A1(\U8/DATA1_17 ), .A2(n374), .ZN(\U7/Z_17 ) );
  AND2_X1 U33 ( .A1(\U8/DATA1_16 ), .A2(n374), .ZN(\U7/Z_16 ) );
  AND2_X1 U34 ( .A1(\U8/DATA1_15 ), .A2(n374), .ZN(\U7/Z_15 ) );
  AND2_X1 U35 ( .A1(\U8/DATA1_14 ), .A2(n374), .ZN(\U7/Z_14 ) );
  OR4_X1 U49 ( .A1(ReadBus[43]), .A2(ReadBus[42]), .A3(ReadBus[45]), .A4(
        ReadBus[44]), .ZN(n22) );
  OAI22_X2 U3 ( .A1(n394), .A2(n440), .B1(n32), .B2(n4), .ZN(n40) );
  OAI22_X2 U5 ( .A1(n2), .A2(n439), .B1(n31), .B2(n4), .ZN(n41) );
  OAI22_X2 U7 ( .A1(n393), .A2(n438), .B1(n30), .B2(n4), .ZN(n42) );
  OAI22_X2 U9 ( .A1(n394), .A2(n437), .B1(n29), .B2(n4), .ZN(n43) );
  OAI22_X2 U11 ( .A1(n2), .A2(n436), .B1(n28), .B2(n4), .ZN(n44) );
  OAI22_X2 U13 ( .A1(n393), .A2(n435), .B1(n27), .B2(n4), .ZN(n45) );
  OAI22_X2 U15 ( .A1(n394), .A2(n434), .B1(n26), .B2(n4), .ZN(n46) );
  OAI22_X2 U19 ( .A1(n2), .A2(\add_63/A[0] ), .B1(n47), .B2(n4), .ZN(n49) );
  NOR3_X2 U43 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n17) );
  NAND3_X2 U44 ( .A1(ReadBus[33]), .A2(ReadBus[31]), .A3(ReadBus[35]), .ZN(n20) );
  NAND3_X2 U45 ( .A1(ReadBus[27]), .A2(ReadBus[25]), .A3(ReadBus[29]), .ZN(n19) );
  NAND4_X2 U46 ( .A1(ReadBus[21]), .A2(start), .A3(ReadBus[23]), .A4(n21), 
        .ZN(n18) );
  NOR4_X2 U47 ( .A1(ReadBus[26]), .A2(ReadBus[24]), .A3(ReadBus[22]), .A4(
        ReadBus[20]), .ZN(n21) );
  NOR4_X2 U48 ( .A1(n22), .A2(ReadBus[39]), .A3(ReadBus[41]), .A4(ReadBus[40]), 
        .ZN(n16) );
  NOR4_X2 U50 ( .A1(ReadBus[38]), .A2(ReadBus[37]), .A3(ReadBus[36]), .A4(
        ReadBus[34]), .ZN(n15) );
  NOR3_X2 U51 ( .A1(ReadBus[28]), .A2(ReadBus[32]), .A3(ReadBus[30]), .ZN(n14)
         );
  DFFR_X2 \ReadAddress_reg[5]  ( .D(\U5/Z_5 ), .CK(clock), .RN(n397), .Q(
        \add_60/A[5] ), .QN(n387) );
  DFFR_X2 \ReadAddress_reg[4]  ( .D(\U5/Z_4 ), .CK(clock), .RN(n396), .Q(
        \add_60/A[4] ), .QN(n386) );
  DFFR_X2 \ReadAddress_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .RN(n396), .Q(
        \add_60/A[2] ), .QN(n384) );
  DFFR_X2 \ReadAddress_reg[0]  ( .D(\U5/Z_0 ), .CK(clock), .RN(n396), .Q(
        \add_60/A[0] ), .QN(n33) );
  DFFR_X2 \ReadAddress_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .RN(n396), .Q(
        \add_60/A[1] ), .QN(n376) );
  DFFR_X2 \ReadAddress_reg[7]  ( .D(\U5/Z_7 ), .CK(clock), .RN(n397), .Q(
        \add_60/A[7] ), .QN(n388) );
  DFFR_X2 \ReadAddress_reg[3]  ( .D(\U5/Z_3 ), .CK(clock), .RN(n396), .Q(
        \add_60/A[3] ), .QN(n385) );
  DFFR_X2 \ReadAddress_reg[9]  ( .D(\U5/Z_9 ), .CK(clock), .RN(n397), .Q(
        \add_60/A[9] ), .QN(n389) );
  DFFR_X2 \count_reg[0]  ( .D(n49), .CK(clock), .RN(n398), .Q(\add_63/A[0] ), 
        .QN(n47) );
  DFFR_X2 \count_reg[4]  ( .D(n43), .CK(clock), .RN(n399), .Q(\add_63/A[4] ), 
        .QN(n29) );
  DFFR_X2 \count_reg[3]  ( .D(n42), .CK(clock), .RN(n399), .Q(\add_63/A[3] ), 
        .QN(n30) );
  DFFR_X2 \count_reg[2]  ( .D(n41), .CK(clock), .RN(n399), .Q(\add_63/A[2] ), 
        .QN(n31) );
  DFFR_X2 \count_reg[1]  ( .D(n40), .CK(clock), .RN(n398), .Q(\add_63/A[1] ), 
        .QN(n32) );
  DFFR_X2 \ReadAddress_reg[11]  ( .D(\U5/Z_11 ), .CK(clock), .RN(n398), .Q(
        \add_60/A[11] ), .QN(n390) );
  DFFR_X2 \count_reg[5]  ( .D(n44), .CK(clock), .RN(n399), .Q(\add_63/A[5] ), 
        .QN(n28) );
  DFFR_X2 \ReadAddress_reg[12]  ( .D(\U5/Z_12 ), .CK(clock), .RN(n398), .Q(
        \add_60/A[12] ), .QN(n391) );
  DFFR_X2 \count_reg[6]  ( .D(n45), .CK(clock), .RN(n399), .Q(\add_63/A[6] ), 
        .QN(n27) );
  DFFR_X2 \count_reg[8]  ( .D(n48), .CK(clock), .RN(n396), .Q(\add_63/A[8] ), 
        .QN(n1) );
  DFFR_X2 \count_reg[7]  ( .D(n46), .CK(clock), .RN(n399), .Q(\add_63/A[7] ), 
        .QN(n26) );
  DFFR_X2 \ReadAddress_reg[13]  ( .D(\U5/Z_13 ), .CK(clock), .RN(n398), .Q(
        \add_60/A[13] ), .QN(n392) );
  DFFR_X2 \ReadAddress_reg[15]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n398), .Q(
        \add_60/A[15] ), .QN(n34) );
  DFFR_X2 done1_reg ( .D(n210), .CK(clock), .RN(reset_n), .Q(n208) );
  DFFR_X2 done_reg ( .D(n208), .CK(clock), .RN(n396), .Q(done) );
  DFFR_X2 \StoreAddress_reg[15]  ( .D(\add_60/A[15] ), .CK(clock), .RN(n398), 
        .Q(StoreAddress[15]) );
  DFFR_X2 \StoreAddress_reg[0]  ( .D(\add_60/A[0] ), .CK(clock), .RN(n396), 
        .Q(StoreAddress[0]) );
  DFFR_X2 \StoreAddress_reg[5]  ( .D(\add_60/A[5] ), .CK(clock), .RN(n397), 
        .Q(StoreAddress[5]) );
  DFFR_X2 \StoreAddress_reg[4]  ( .D(\add_60/A[4] ), .CK(clock), .RN(n396), 
        .Q(StoreAddress[4]) );
  DFFR_X2 \StoreAddress_reg[2]  ( .D(\add_60/A[2] ), .CK(clock), .RN(n396), 
        .Q(StoreAddress[2]) );
  DFFR_X2 \StoreAddress_reg[1]  ( .D(\add_60/A[1] ), .CK(clock), .RN(n396), 
        .Q(StoreAddress[1]) );
  DFFR_X2 \StoreAddress_reg[13]  ( .D(\add_60/A[13] ), .CK(clock), .RN(n398), 
        .Q(StoreAddress[13]) );
  DFFR_X2 \StoreAddress_reg[12]  ( .D(\add_60/A[12] ), .CK(clock), .RN(n398), 
        .Q(StoreAddress[12]) );
  DFFR_X2 \StoreAddress_reg[11]  ( .D(\add_60/A[11] ), .CK(clock), .RN(n398), 
        .Q(StoreAddress[11]) );
  DFFR_X2 \StoreAddress_reg[9]  ( .D(\add_60/A[9] ), .CK(clock), .RN(n397), 
        .Q(StoreAddress[9]) );
  DFFR_X2 \StoreAddress_reg[7]  ( .D(\add_60/A[7] ), .CK(clock), .RN(n397), 
        .Q(StoreAddress[7]) );
  DFFR_X2 \StoreAddress_reg[3]  ( .D(\add_60/A[3] ), .CK(clock), .RN(n396), 
        .Q(StoreAddress[3]) );
  DFFR_X2 \StoreAddress_reg[10]  ( .D(\add_60/A[10] ), .CK(clock), .RN(n397), 
        .Q(StoreAddress[10]) );
  DFFR_X2 \StoreAddress_reg[8]  ( .D(\add_60/A[8] ), .CK(clock), .RN(n397), 
        .Q(StoreAddress[8]) );
  DFFR_X2 \StoreAddress_reg[6]  ( .D(\add_60/A[6] ), .CK(clock), .RN(n397), 
        .Q(StoreAddress[6]) );
  DFFR_X2 \StoreAddress_reg[14]  ( .D(\add_60/A[14] ), .CK(clock), .RN(n398), 
        .Q(StoreAddress[14]) );
  DFFR_X2 \ReadAddress_reg[6]  ( .D(\U5/Z_6 ), .CK(clock), .RN(n397), .Q(
        \add_60/A[6] ) );
  DFFR_X2 \ReadAddress_reg[8]  ( .D(\U5/Z_8 ), .CK(clock), .RN(n397), .Q(
        \add_60/A[8] ) );
  DFFR_X2 \AccumlateOut_reg[19]  ( .D(\U7/Z_19 ), .CK(clock), .RN(n399), .Q(
        AccumlateOut[19]) );
  DFFR_X2 \AccumlateOut_reg[18]  ( .D(\U7/Z_18 ), .CK(clock), .RN(n399), .Q(
        AccumlateOut[18]) );
  DFFR_X2 \AccumlateOut_reg[17]  ( .D(\U7/Z_17 ), .CK(clock), .RN(n399), .Q(
        AccumlateOut[17]) );
  DFFR_X2 \AccumlateOut_reg[16]  ( .D(\U7/Z_16 ), .CK(clock), .RN(n399), .Q(
        AccumlateOut[16]) );
  DFFR_X2 \AccumlateOut_reg[15]  ( .D(\U7/Z_15 ), .CK(clock), .RN(n399), .Q(
        AccumlateOut[15]) );
  DFFR_X2 \AccumlateOut_reg[14]  ( .D(\U7/Z_14 ), .CK(clock), .RN(n399), .Q(
        AccumlateOut[14]) );
  DFFR_X2 \AccumlateOut_reg[13]  ( .D(\U7/Z_13 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[13]) );
  DFFR_X2 \AccumlateOut_reg[12]  ( .D(\U7/Z_12 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[12]) );
  DFFR_X2 \AccumlateOut_reg[11]  ( .D(\U7/Z_11 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[11]) );
  DFFR_X2 \AccumlateOut_reg[10]  ( .D(\U7/Z_10 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[10]) );
  DFFR_X2 \AccumlateOut_reg[9]  ( .D(\U7/Z_9 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[9]) );
  DFFR_X2 \AccumlateOut_reg[8]  ( .D(\U7/Z_8 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[8]) );
  DFFR_X2 \AccumlateOut_reg[7]  ( .D(\U7/Z_7 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[7]) );
  DFFR_X2 \AccumlateOut_reg[6]  ( .D(\U7/Z_6 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[6]) );
  DFFR_X2 \AccumlateOut_reg[5]  ( .D(\U7/Z_5 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[5]) );
  DFFR_X2 \AccumlateOut_reg[3]  ( .D(\U7/Z_3 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[3]) );
  DFFR_X2 \AccumlateOut_reg[2]  ( .D(\U7/Z_2 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[2]) );
  DFFR_X2 \ReadAddress_reg[14]  ( .D(\U5/Z_14 ), .CK(clock), .RN(n398), .Q(
        \add_60/A[14] ), .QN(n428) );
  DFFR_X2 \ReadAddress_reg[10]  ( .D(\U5/Z_10 ), .CK(clock), .RN(n397), .Q(
        \add_60/A[10] ) );
  DFFR_X2 \AccumlateOut_reg[4]  ( .D(\U7/Z_4 ), .CK(clock), .RN(n400), .Q(
        AccumlateOut[4]) );
  DFFR_X2 \AccumlateOut_reg[1]  ( .D(\U7/Z_1 ), .CK(clock), .RN(reset_n), .Q(
        AccumlateOut[1]) );
  DFFR_X2 \AccumlateOut_reg[0]  ( .D(\U7/Z_0 ), .CK(clock), .RN(reset_n), .Q(
        AccumlateOut[0]) );
  AND4_X4 U4 ( .A1(n16), .A2(n17), .A3(n14), .A4(n15), .ZN(n374) );
  NOR2_X2 U6 ( .A1(n429), .A2(n428), .ZN(n430) );
  OR2_X4 U8 ( .A1(n392), .A2(n426), .ZN(n429) );
  INV_X2 U10 ( .A(n416), .ZN(n379) );
  NAND2_X2 U12 ( .A1(\add_60/A[8] ), .A2(n379), .ZN(n418) );
  NAND2_X2 U14 ( .A1(n375), .A2(n380), .ZN(n408) );
  OR2_X4 U16 ( .A1(n390), .A2(n422), .ZN(n424) );
  INV_X1 U17 ( .A(n375), .ZN(n404) );
  NOR2_X2 U18 ( .A1(n376), .A2(n33), .ZN(n375) );
  NOR2_X2 U20 ( .A1(n389), .A2(n418), .ZN(n377) );
  NOR2_X2 U21 ( .A1(n387), .A2(n410), .ZN(n378) );
  OR2_X4 U22 ( .A1(n386), .A2(n408), .ZN(n410) );
  NAND2_X2 U23 ( .A1(\add_60/A[6] ), .A2(n378), .ZN(n414) );
  NAND2_X2 U24 ( .A1(\add_60/A[10] ), .A2(n377), .ZN(n422) );
  NOR2_X2 U25 ( .A1(n384), .A2(n385), .ZN(n380) );
  NAND2_X2 U26 ( .A1(n34), .A2(n381), .ZN(n382) );
  NAND2_X1 U27 ( .A1(\add_60/A[15] ), .A2(n430), .ZN(n383) );
  NAND2_X2 U28 ( .A1(n382), .A2(n383), .ZN(n432) );
  INV_X2 U29 ( .A(n430), .ZN(n381) );
  INV_X4 U36 ( .A(n401), .ZN(n400) );
  INV_X4 U37 ( .A(n401), .ZN(n399) );
  INV_X4 U38 ( .A(n401), .ZN(n397) );
  INV_X4 U39 ( .A(n401), .ZN(n396) );
  INV_X4 U40 ( .A(n401), .ZN(n398) );
  INV_X4 U41 ( .A(reset_n), .ZN(n401) );
  INV_X4 U42 ( .A(start), .ZN(n395) );
  NAND2_X2 U52 ( .A1(n393), .A2(start), .ZN(n4) );
  OAI21_X2 U53 ( .B1(n433), .B2(n394), .A(n4), .ZN(n48) );
  OR2_X1 U54 ( .A1(n384), .A2(n404), .ZN(n406) );
  OR2_X1 U55 ( .A1(n387), .A2(n410), .ZN(n412) );
  OR2_X1 U56 ( .A1(n388), .A2(n414), .ZN(n416) );
  OR2_X1 U57 ( .A1(n389), .A2(n418), .ZN(n420) );
  OR2_X1 U58 ( .A1(n391), .A2(n424), .ZN(n426) );
  NAND2_X2 U59 ( .A1(start), .A2(n1), .ZN(n393) );
  NAND2_X2 U60 ( .A1(start), .A2(n1), .ZN(n394) );
  NAND2_X2 U61 ( .A1(start), .A2(n1), .ZN(n2) );
  INV_X4 U62 ( .A(\U3/U1/DATA1_7 ), .ZN(n434) );
  INV_X4 U63 ( .A(\U3/U1/DATA1_6 ), .ZN(n435) );
  INV_X4 U64 ( .A(\U3/U1/DATA1_5 ), .ZN(n436) );
  INV_X4 U65 ( .A(\U3/U1/DATA1_4 ), .ZN(n437) );
  INV_X4 U66 ( .A(\U3/U1/DATA1_3 ), .ZN(n438) );
  INV_X4 U67 ( .A(\U3/U1/DATA1_2 ), .ZN(n439) );
  INV_X4 U68 ( .A(\U3/U1/DATA1_1 ), .ZN(n440) );
  NOR2_X2 U69 ( .A1(\add_60/A[0] ), .A2(n2), .ZN(\U5/Z_0 ) );
  XNOR2_X2 U70 ( .A(\add_60/A[0] ), .B(\add_60/A[1] ), .ZN(n402) );
  NOR2_X2 U71 ( .A1(n393), .A2(n402), .ZN(\U5/Z_1 ) );
  XOR2_X2 U72 ( .A(n404), .B(\add_60/A[2] ), .Z(n403) );
  NOR2_X2 U73 ( .A1(n2), .A2(n403), .ZN(\U5/Z_2 ) );
  XOR2_X2 U74 ( .A(n406), .B(\add_60/A[3] ), .Z(n405) );
  NOR2_X2 U77 ( .A1(n2), .A2(n405), .ZN(\U5/Z_3 ) );
  XOR2_X2 U78 ( .A(n408), .B(\add_60/A[4] ), .Z(n407) );
  NOR2_X2 U79 ( .A1(n393), .A2(n407), .ZN(\U5/Z_4 ) );
  XOR2_X2 U80 ( .A(n410), .B(\add_60/A[5] ), .Z(n409) );
  NOR2_X2 U81 ( .A1(n394), .A2(n409), .ZN(\U5/Z_5 ) );
  XOR2_X2 U82 ( .A(n412), .B(\add_60/A[6] ), .Z(n411) );
  NOR2_X2 U83 ( .A1(n2), .A2(n411), .ZN(\U5/Z_6 ) );
  XOR2_X2 U84 ( .A(n414), .B(\add_60/A[7] ), .Z(n413) );
  NOR2_X2 U85 ( .A1(n393), .A2(n413), .ZN(\U5/Z_7 ) );
  XOR2_X2 U86 ( .A(n416), .B(\add_60/A[8] ), .Z(n415) );
  NOR2_X2 U87 ( .A1(n394), .A2(n415), .ZN(\U5/Z_8 ) );
  XOR2_X2 U88 ( .A(n418), .B(\add_60/A[9] ), .Z(n417) );
  NOR2_X2 U89 ( .A1(n2), .A2(n417), .ZN(\U5/Z_9 ) );
  XOR2_X2 U90 ( .A(n420), .B(\add_60/A[10] ), .Z(n419) );
  NOR2_X2 U91 ( .A1(n393), .A2(n419), .ZN(\U5/Z_10 ) );
  XOR2_X2 U92 ( .A(n422), .B(\add_60/A[11] ), .Z(n421) );
  NOR2_X2 U93 ( .A1(n394), .A2(n421), .ZN(\U5/Z_11 ) );
  XOR2_X2 U94 ( .A(n424), .B(\add_60/A[12] ), .Z(n423) );
  NOR2_X2 U95 ( .A1(n2), .A2(n423), .ZN(\U5/Z_12 ) );
  XOR2_X2 U96 ( .A(n426), .B(\add_60/A[13] ), .Z(n425) );
  NOR2_X2 U97 ( .A1(n393), .A2(n425), .ZN(\U5/Z_13 ) );
  XOR2_X2 U98 ( .A(n429), .B(\add_60/A[14] ), .Z(n427) );
  NOR2_X2 U99 ( .A1(n394), .A2(n427), .ZN(\U5/Z_14 ) );
  INV_X4 U100 ( .A(\U4/DATA3_0 ), .ZN(n431) );
  OAI22_X2 U101 ( .A1(n393), .A2(n432), .B1(start), .B2(n431), .ZN(\U4/Z_0 )
         );
  AND2_X1 U102 ( .A1(\U8/DATA1_0 ), .A2(n374), .ZN(\U7/Z_0 ) );
  AND2_X1 U103 ( .A1(\U8/DATA1_1 ), .A2(n374), .ZN(\U7/Z_1 ) );
  AND2_X1 U104 ( .A1(\U8/DATA1_2 ), .A2(n374), .ZN(\U7/Z_2 ) );
  AND2_X1 U105 ( .A1(\U8/DATA1_3 ), .A2(n374), .ZN(\U7/Z_3 ) );
  AND2_X1 U106 ( .A1(\U8/DATA1_4 ), .A2(n374), .ZN(\U7/Z_4 ) );
  AND2_X1 U107 ( .A1(\U8/DATA1_5 ), .A2(n374), .ZN(\U7/Z_5 ) );
  AND2_X1 U108 ( .A1(\U8/DATA1_6 ), .A2(n374), .ZN(\U7/Z_6 ) );
  AND2_X1 U109 ( .A1(\U8/DATA1_7 ), .A2(n374), .ZN(\U7/Z_7 ) );
  AND2_X1 U110 ( .A1(\U8/DATA1_8 ), .A2(n374), .ZN(\U7/Z_8 ) );
  AND2_X1 U111 ( .A1(\U8/DATA1_9 ), .A2(n374), .ZN(\U7/Z_9 ) );
  AND2_X1 U112 ( .A1(\U8/DATA1_10 ), .A2(n374), .ZN(\U7/Z_10 ) );
  AND2_X1 U113 ( .A1(\U8/DATA1_11 ), .A2(n374), .ZN(\U7/Z_11 ) );
  AND2_X1 U114 ( .A1(\U8/DATA1_12 ), .A2(n374), .ZN(\U7/Z_12 ) );
  AND2_X1 U115 ( .A1(\U8/DATA1_13 ), .A2(n374), .ZN(\U7/Z_13 ) );
  INV_X4 U116 ( .A(\add_63/carry[8] ), .ZN(n433) );
endmodule


module Cdf_Accumlate ( clock, reset_n, AccumlateIn, StartIn, StoreAddressIn, 
        AccumlateResult, StoreAddressOut, StartOut, CdfMin, CdfValid );
  input [19:0] AccumlateIn;
  input [15:0] StoreAddressIn;
  output [19:0] AccumlateResult;
  output [15:0] StoreAddressOut;
  output [19:0] CdfMin;
  input clock, reset_n, StartIn;
  output StartOut, CdfValid;
  wire   \U10/DATA2_0 , \U10/DATA2_1 , \U10/DATA2_2 , \U10/DATA2_3 ,
         \U10/DATA2_4 , \U10/DATA2_5 , \U10/DATA2_6 , \U10/DATA2_7 ,
         \U10/DATA2_8 , \U10/DATA2_9 , \U10/DATA2_10 , \U10/DATA2_11 ,
         \U10/DATA2_12 , \U10/DATA2_13 , \U10/DATA2_14 , \U10/DATA2_15 ,
         \U10/DATA2_16 , \U10/DATA2_17 , \U10/DATA2_18 , \U10/DATA2_19 ,
         \U10/DATA1_0 , \U10/DATA1_1 , \U10/DATA1_2 , \U10/DATA1_3 ,
         \U10/DATA1_4 , \U10/DATA1_5 , \U10/DATA1_6 , \U10/DATA1_7 ,
         \U10/DATA1_8 , \U10/DATA1_9 , \U10/DATA1_10 , \U10/DATA1_11 ,
         \U10/DATA1_12 , \U10/DATA1_13 , \U10/DATA1_14 , \U10/DATA1_15 ,
         \U10/DATA1_16 , \U10/DATA1_17 , \U10/DATA1_18 , \U10/DATA1_19 ,
         \U8/Z_0 , \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 ,
         \U4/Z_6 , \U4/Z_7 , \U4/Z_8 , \U4/Z_9 , \U4/Z_10 , \U4/Z_11 ,
         \U4/Z_12 , \U4/Z_13 , \U4/Z_14 , \U4/Z_15 , \U4/Z_16 , \U4/Z_17 ,
         \U4/Z_18 , \U4/Z_19 , \add_48/B[0] , \add_48/B[1] , \add_48/B[2] ,
         \add_48/B[3] , \add_48/B[4] , \add_48/B[5] , \add_48/B[6] ,
         \add_48/B[7] , \add_48/B[8] , \add_48/B[9] , \add_48/B[10] ,
         \add_48/B[11] , \add_48/B[12] , \add_48/B[13] , \add_48/B[14] ,
         \add_48/B[15] , \add_48/B[16] , \add_48/B[17] , \add_48/B[18] ,
         \add_48/B[19] , n5, n6, n11, n16, n17, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n43, n44, n45, n48, n49, n50, n51, n52, n53, n54, n55, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n217, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391;
  assign CdfMin[0] = \U10/DATA2_0 ;
  assign CdfMin[1] = \U10/DATA2_1 ;
  assign CdfMin[2] = \U10/DATA2_2 ;
  assign CdfMin[3] = \U10/DATA2_3 ;
  assign CdfMin[4] = \U10/DATA2_4 ;
  assign CdfMin[5] = \U10/DATA2_5 ;
  assign CdfMin[6] = \U10/DATA2_6 ;
  assign CdfMin[7] = \U10/DATA2_7 ;
  assign CdfMin[8] = \U10/DATA2_8 ;
  assign CdfMin[9] = \U10/DATA2_9 ;
  assign CdfMin[10] = \U10/DATA2_10 ;
  assign CdfMin[11] = \U10/DATA2_11 ;
  assign CdfMin[12] = \U10/DATA2_12 ;
  assign CdfMin[13] = \U10/DATA2_13 ;
  assign CdfMin[14] = \U10/DATA2_14 ;
  assign CdfMin[15] = \U10/DATA2_15 ;
  assign CdfMin[16] = \U10/DATA2_16 ;
  assign CdfMin[17] = \U10/DATA2_17 ;
  assign CdfMin[18] = \U10/DATA2_18 ;
  assign CdfMin[19] = \U10/DATA2_19 ;
  assign AccumlateResult[0] = \U10/DATA1_0 ;
  assign AccumlateResult[1] = \U10/DATA1_1 ;
  assign AccumlateResult[2] = \U10/DATA1_2 ;
  assign AccumlateResult[3] = \U10/DATA1_3 ;
  assign AccumlateResult[4] = \U10/DATA1_4 ;
  assign AccumlateResult[5] = \U10/DATA1_5 ;
  assign AccumlateResult[6] = \U10/DATA1_6 ;
  assign AccumlateResult[7] = \U10/DATA1_7 ;
  assign AccumlateResult[8] = \U10/DATA1_8 ;
  assign AccumlateResult[9] = \U10/DATA1_9 ;
  assign AccumlateResult[10] = \U10/DATA1_10 ;
  assign AccumlateResult[11] = \U10/DATA1_11 ;
  assign AccumlateResult[12] = \U10/DATA1_12 ;
  assign AccumlateResult[13] = \U10/DATA1_13 ;
  assign AccumlateResult[14] = \U10/DATA1_14 ;
  assign AccumlateResult[15] = \U10/DATA1_15 ;
  assign AccumlateResult[16] = \U10/DATA1_16 ;
  assign AccumlateResult[17] = \U10/DATA1_17 ;
  assign AccumlateResult[18] = \U10/DATA1_18 ;
  assign AccumlateResult[19] = \U10/DATA1_19 ;
  assign \add_48/B[0]  = AccumlateIn[0];
  assign \add_48/B[1]  = AccumlateIn[1];
  assign \add_48/B[2]  = AccumlateIn[2];
  assign \add_48/B[3]  = AccumlateIn[3];
  assign \add_48/B[4]  = AccumlateIn[4];
  assign \add_48/B[5]  = AccumlateIn[5];
  assign \add_48/B[6]  = AccumlateIn[6];
  assign \add_48/B[7]  = AccumlateIn[7];
  assign \add_48/B[8]  = AccumlateIn[8];
  assign \add_48/B[9]  = AccumlateIn[9];
  assign \add_48/B[10]  = AccumlateIn[10];
  assign \add_48/B[11]  = AccumlateIn[11];
  assign \add_48/B[12]  = AccumlateIn[12];
  assign \add_48/B[13]  = AccumlateIn[13];
  assign \add_48/B[14]  = AccumlateIn[14];
  assign \add_48/B[15]  = AccumlateIn[15];
  assign \add_48/B[16]  = AccumlateIn[16];
  assign \add_48/B[17]  = AccumlateIn[17];
  assign \add_48/B[18]  = AccumlateIn[18];
  assign \add_48/B[19]  = AccumlateIn[19];

  DFF_X1 \StoreAddressOut_reg[15]  ( .D(StoreAddressIn[15]), .CK(clock), .Q(
        StoreAddressOut[15]) );
  DFF_X1 \StoreAddressOut_reg[14]  ( .D(StoreAddressIn[14]), .CK(clock), .Q(
        StoreAddressOut[14]) );
  DFF_X1 \StoreAddressOut_reg[13]  ( .D(StoreAddressIn[13]), .CK(clock), .Q(
        StoreAddressOut[13]) );
  DFF_X1 \StoreAddressOut_reg[12]  ( .D(StoreAddressIn[12]), .CK(clock), .Q(
        StoreAddressOut[12]) );
  DFF_X1 \StoreAddressOut_reg[11]  ( .D(StoreAddressIn[11]), .CK(clock), .Q(
        StoreAddressOut[11]) );
  DFF_X1 \StoreAddressOut_reg[10]  ( .D(StoreAddressIn[10]), .CK(clock), .Q(
        StoreAddressOut[10]) );
  DFF_X1 \StoreAddressOut_reg[9]  ( .D(StoreAddressIn[9]), .CK(clock), .Q(
        StoreAddressOut[9]) );
  DFF_X1 \StoreAddressOut_reg[8]  ( .D(StoreAddressIn[8]), .CK(clock), .Q(
        StoreAddressOut[8]) );
  DFF_X1 \StoreAddressOut_reg[7]  ( .D(StoreAddressIn[7]), .CK(clock), .Q(
        StoreAddressOut[7]) );
  DFF_X1 \StoreAddressOut_reg[6]  ( .D(StoreAddressIn[6]), .CK(clock), .Q(
        StoreAddressOut[6]) );
  DFF_X1 \StoreAddressOut_reg[5]  ( .D(StoreAddressIn[5]), .CK(clock), .Q(
        StoreAddressOut[5]) );
  DFF_X1 \StoreAddressOut_reg[4]  ( .D(StoreAddressIn[4]), .CK(clock), .Q(
        StoreAddressOut[4]) );
  DFF_X1 \StoreAddressOut_reg[3]  ( .D(StoreAddressIn[3]), .CK(clock), .Q(
        StoreAddressOut[3]) );
  DFF_X1 \StoreAddressOut_reg[2]  ( .D(StoreAddressIn[2]), .CK(clock), .Q(
        StoreAddressOut[2]) );
  DFF_X1 \StoreAddressOut_reg[1]  ( .D(StoreAddressIn[1]), .CK(clock), .Q(
        StoreAddressOut[1]) );
  DFF_X1 \StoreAddressOut_reg[0]  ( .D(StoreAddressIn[0]), .CK(clock), .Q(
        StoreAddressOut[0]) );
  NAND2_X2 U24 ( .A1(StartIn), .A2(n43), .ZN(n44) );
  NAND4_X2 U27 ( .A1(n48), .A2(n49), .A3(n50), .A4(n51), .ZN(n45) );
  NOR3_X2 U28 ( .A1(n52), .A2(\U10/DATA2_6 ), .A3(\U10/DATA2_5 ), .ZN(n51) );
  NAND3_X2 U29 ( .A1(n33), .A2(n32), .A3(n34), .ZN(n52) );
  NOR3_X2 U30 ( .A1(n53), .A2(\U10/DATA2_19 ), .A3(\U10/DATA2_18 ), .ZN(n50)
         );
  NAND3_X2 U31 ( .A1(n38), .A2(n37), .A3(n39), .ZN(n53) );
  NOR3_X2 U32 ( .A1(n54), .A2(\U10/DATA2_14 ), .A3(\U10/DATA2_13 ), .ZN(n49)
         );
  NAND3_X2 U33 ( .A1(n25), .A2(n24), .A3(n26), .ZN(n54) );
  NOR3_X2 U34 ( .A1(n55), .A2(\U10/DATA2_1 ), .A3(\U10/DATA2_0 ), .ZN(n48) );
  NAND3_X2 U35 ( .A1(n30), .A2(n29), .A3(n31), .ZN(n55) );
  DFFR_X2 \AccumlateResult_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .RN(reset_n), 
        .Q(\U10/DATA1_0 ), .QN(n21) );
  DFFR_X2 \AccumlateResult_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .RN(reset_n), 
        .Q(\U10/DATA1_1 ), .QN(n20) );
  DFFR_X2 \AccumlateResult_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(reset_n), 
        .Q(\U10/DATA1_4 ), .QN(n17) );
  DFFR_X2 \AccumlateResult_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n244), .Q(
        \U10/DATA1_5 ), .QN(n16) );
  DFFR_X2 \AccumlateResult_reg[18]  ( .D(\U4/Z_18 ), .CK(clock), .RN(n243), 
        .Q(\U10/DATA1_18 ), .QN(n379) );
  DFFR_X2 \AccumlateResult_reg[17]  ( .D(\U4/Z_17 ), .CK(clock), .RN(n243), 
        .Q(\U10/DATA1_17 ), .QN(n380) );
  DFFR_X2 \AccumlateResult_reg[19]  ( .D(\U4/Z_19 ), .CK(clock), .RN(n243), 
        .Q(\U10/DATA1_19 ), .QN(n366) );
  DFFR_X2 \AccumlateResult_reg[16]  ( .D(\U4/Z_16 ), .CK(clock), .RN(n244), 
        .Q(\U10/DATA1_16 ), .QN(n5) );
  DFFR_X2 \AccumlateResult_reg[15]  ( .D(\U4/Z_15 ), .CK(clock), .RN(n244), 
        .Q(\U10/DATA1_15 ), .QN(n6) );
  DFFR_X2 \AccumlateResult_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .RN(reset_n), 
        .Q(\U10/DATA1_2 ), .QN(n256) );
  DFFR_X2 \AccumlateResult_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(reset_n), 
        .Q(\U10/DATA1_3 ), .QN(n262) );
  DFFR_X2 \AccumlateResult_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n244), .Q(
        \U10/DATA1_6 ), .QN(n290) );
  DFFR_X2 \CdfMin_reg[14]  ( .D(n67), .CK(clock), .RN(n243), .Q(\U10/DATA2_14 ), .QN(n27) );
  DFFR_X2 \CdfMin_reg[2]  ( .D(n79), .CK(clock), .RN(n242), .Q(\U10/DATA2_2 ), 
        .QN(n39) );
  DFFR_X2 \CdfMin_reg[11]  ( .D(n70), .CK(clock), .RN(n242), .Q(\U10/DATA2_11 ), .QN(n30) );
  DFFR_X2 \CdfMin_reg[17]  ( .D(n64), .CK(clock), .RN(n243), .Q(\U10/DATA2_17 ), .QN(n24) );
  DFFR_X2 \CdfMin_reg[8]  ( .D(n73), .CK(clock), .RN(n242), .Q(\U10/DATA2_8 ), 
        .QN(n33) );
  DFFR_X2 \CdfMin_reg[5]  ( .D(n76), .CK(clock), .RN(n242), .Q(\U10/DATA2_5 ), 
        .QN(n36) );
  DFFR_X2 \CdfMin_reg[13]  ( .D(n68), .CK(clock), .RN(n243), .Q(\U10/DATA2_13 ), .QN(n28) );
  DFFR_X2 \CdfMin_reg[10]  ( .D(n71), .CK(clock), .RN(n242), .Q(\U10/DATA2_10 ), .QN(n31) );
  DFFR_X2 \CdfMin_reg[12]  ( .D(n69), .CK(clock), .RN(n243), .Q(\U10/DATA2_12 ), .QN(n29) );
  DFFR_X2 \CdfMin_reg[3]  ( .D(n78), .CK(clock), .RN(n242), .Q(\U10/DATA2_3 ), 
        .QN(n38) );
  DFFR_X2 \CdfMin_reg[9]  ( .D(n72), .CK(clock), .RN(n242), .Q(\U10/DATA2_9 ), 
        .QN(n32) );
  DFFR_X2 \CdfMin_reg[6]  ( .D(n75), .CK(clock), .RN(n242), .Q(\U10/DATA2_6 ), 
        .QN(n35) );
  DFFR_X2 \CdfMin_reg[18]  ( .D(n63), .CK(clock), .RN(n243), .Q(\U10/DATA2_18 ), .QN(n23) );
  DFFR_X2 \CdfMin_reg[7]  ( .D(n74), .CK(clock), .RN(n242), .Q(\U10/DATA2_7 ), 
        .QN(n34) );
  DFFR_X2 \CdfMin_reg[16]  ( .D(n65), .CK(clock), .RN(n243), .Q(\U10/DATA2_16 ), .QN(n25) );
  DFFR_X2 \CdfMin_reg[1]  ( .D(n80), .CK(clock), .RN(n242), .Q(\U10/DATA2_1 ), 
        .QN(n40) );
  DFFR_X2 \CdfMin_reg[19]  ( .D(n62), .CK(clock), .RN(n243), .Q(\U10/DATA2_19 ), .QN(n22) );
  DFFR_X2 \CdfMin_reg[15]  ( .D(n66), .CK(clock), .RN(n243), .Q(\U10/DATA2_15 ), .QN(n26) );
  DFFR_X2 \CdfMin_reg[4]  ( .D(n77), .CK(clock), .RN(n242), .Q(\U10/DATA2_4 ), 
        .QN(n37) );
  DFFR_X2 \CdfMin_reg[0]  ( .D(n81), .CK(clock), .RN(n243), .Q(\U10/DATA2_0 ), 
        .QN(n41) );
  DFFR_X2 \AccumlateResult_reg[8]  ( .D(\U4/Z_8 ), .CK(clock), .RN(n244), .Q(
        \U10/DATA1_8 ), .QN(n385) );
  DFFR_X2 \AccumlateResult_reg[7]  ( .D(\U4/Z_7 ), .CK(clock), .RN(n244), .Q(
        \U10/DATA1_7 ), .QN(n298) );
  DFFR_X2 \AccumlateResult_reg[9]  ( .D(\U4/Z_9 ), .CK(clock), .RN(n244), .Q(
        \U10/DATA1_9 ), .QN(n384) );
  DFFR_X2 \AccumlateResult_reg[10]  ( .D(\U4/Z_10 ), .CK(clock), .RN(n244), 
        .Q(\U10/DATA1_10 ), .QN(n11) );
  DFFR_X2 \AccumlateResult_reg[11]  ( .D(\U4/Z_11 ), .CK(clock), .RN(n244), 
        .Q(\U10/DATA1_11 ), .QN(n323) );
  DFFR_X2 \AccumlateResult_reg[12]  ( .D(\U4/Z_12 ), .CK(clock), .RN(n244), 
        .Q(\U10/DATA1_12 ), .QN(n329) );
  DFFR_X2 \AccumlateResult_reg[13]  ( .D(\U4/Z_13 ), .CK(clock), .RN(n244), 
        .Q(\U10/DATA1_13 ), .QN(n336) );
  DFFR_X2 \AccumlateResult_reg[14]  ( .D(\U4/Z_14 ), .CK(clock), .RN(n244), 
        .Q(\U10/DATA1_14 ), .QN(n341) );
  DFFR_X2 StartOut_reg ( .D(StartIn), .CK(clock), .RN(reset_n), .Q(StartOut)
         );
  DFFR_X2 CdfValid_reg ( .D(\U8/Z_0 ), .CK(clock), .RN(n242), .Q(CdfValid) );
  AOI22_X4 U3 ( .A1(n332), .A2(n331), .B1(\U10/DATA1_12 ), .B2(\add_48/B[12] ), 
        .ZN(n337) );
  OAI21_X2 U4 ( .B1(\add_48/B[5] ), .B2(\U10/DATA1_5 ), .A(n275), .ZN(n276) );
  INV_X4 U5 ( .A(\add_48/B[10] ), .ZN(n222) );
  AOI22_X2 U6 ( .A1(n349), .A2(n348), .B1(\U10/DATA1_15 ), .B2(\add_48/B[15] ), 
        .ZN(n354) );
  NOR3_X2 U7 ( .A1(n364), .A2(n363), .A3(n362), .ZN(\U4/Z_18 ) );
  OAI211_X4 U8 ( .C1(n301), .C2(n302), .A(n300), .B(n299), .ZN(n311) );
  AND3_X4 U9 ( .A1(n358), .A2(n369), .A3(n361), .ZN(n217) );
  OAI22_X2 U10 ( .A1(n223), .A2(n221), .B1(n11), .B2(n222), .ZN(n220) );
  INV_X1 U11 ( .A(n220), .ZN(n324) );
  INV_X1 U12 ( .A(n224), .ZN(n342) );
  INV_X4 U13 ( .A(n319), .ZN(n221) );
  NOR2_X2 U14 ( .A1(\U10/DATA1_10 ), .A2(\add_48/B[10] ), .ZN(n223) );
  OAI22_X2 U15 ( .A1(n225), .A2(n337), .B1(n336), .B2(n335), .ZN(n224) );
  AND2_X4 U16 ( .A1(n336), .A2(n335), .ZN(n225) );
  AOI221_X2 U17 ( .B1(n233), .B2(n384), .C1(n311), .C2(n235), .A(n234), .ZN(
        n232) );
  NOR2_X1 U18 ( .A1(n361), .A2(n368), .ZN(n226) );
  NOR2_X2 U19 ( .A1(n360), .A2(n359), .ZN(n227) );
  OR3_X2 U20 ( .A1(n226), .A2(n227), .A3(n217), .ZN(n364) );
  INV_X1 U21 ( .A(n361), .ZN(n360) );
  INV_X4 U22 ( .A(n314), .ZN(n234) );
  INV_X4 U23 ( .A(n232), .ZN(n315) );
  INV_X4 U25 ( .A(\add_48/B[9] ), .ZN(n233) );
  OAI221_X2 U26 ( .B1(n373), .B2(n372), .C1(n371), .C2(n370), .A(StartIn), 
        .ZN(n374) );
  XNOR2_X1 U36 ( .A(n358), .B(n236), .ZN(n355) );
  XOR2_X1 U37 ( .A(\add_48/B[8] ), .B(\U10/DATA1_8 ), .Z(n303) );
  XNOR2_X2 U38 ( .A(n228), .B(n293), .ZN(n294) );
  XOR2_X1 U39 ( .A(\add_48/B[7] ), .B(\U10/DATA1_7 ), .Z(n228) );
  XOR2_X1 U40 ( .A(\add_48/B[6] ), .B(\U10/DATA1_6 ), .Z(n287) );
  XOR2_X1 U41 ( .A(\add_48/B[2] ), .B(\U10/DATA1_2 ), .Z(n253) );
  XNOR2_X2 U42 ( .A(n229), .B(n259), .ZN(n260) );
  XOR2_X1 U43 ( .A(\add_48/B[3] ), .B(\U10/DATA1_3 ), .Z(n229) );
  AND2_X4 U44 ( .A1(n377), .A2(n378), .ZN(n230) );
  AND2_X4 U45 ( .A1(n376), .A2(n375), .ZN(n231) );
  NOR3_X2 U46 ( .A1(n230), .A2(n231), .A3(n374), .ZN(\U4/Z_19 ) );
  INV_X4 U47 ( .A(n377), .ZN(n376) );
  INV_X2 U48 ( .A(n373), .ZN(n375) );
  AND2_X4 U49 ( .A1(n313), .A2(n312), .ZN(n235) );
  INV_X4 U50 ( .A(n245), .ZN(n243) );
  INV_X4 U51 ( .A(n245), .ZN(n244) );
  INV_X4 U52 ( .A(n245), .ZN(n242) );
  INV_X4 U53 ( .A(reset_n), .ZN(n245) );
  XNOR2_X2 U54 ( .A(\add_48/B[17] ), .B(\U10/DATA1_17 ), .ZN(n236) );
  NAND2_X2 U55 ( .A1(n251), .A2(n252), .ZN(n263) );
  NAND2_X2 U56 ( .A1(StartIn), .A2(n45), .ZN(n239) );
  NAND2_X2 U57 ( .A1(StartIn), .A2(n45), .ZN(n238) );
  NAND2_X2 U58 ( .A1(StartIn), .A2(n45), .ZN(n43) );
  XNOR2_X2 U59 ( .A(n306), .B(n303), .ZN(n304) );
  XNOR2_X2 U60 ( .A(n270), .B(n267), .ZN(n268) );
  XNOR2_X2 U61 ( .A(n291), .B(n287), .ZN(n288) );
  INV_X4 U62 ( .A(StartIn), .ZN(n362) );
  XNOR2_X2 U63 ( .A(n257), .B(n253), .ZN(n254) );
  XOR2_X1 U64 ( .A(\add_48/B[4] ), .B(\U10/DATA1_4 ), .Z(n267) );
  NAND2_X1 U65 ( .A1(\add_48/B[4] ), .A2(\U10/DATA1_4 ), .ZN(n281) );
  NAND2_X2 U66 ( .A1(\add_48/B[1] ), .A2(\U10/DATA1_1 ), .ZN(n264) );
  XOR2_X1 U67 ( .A(n337), .B(n333), .Z(n334) );
  INV_X2 U68 ( .A(n21), .ZN(n237) );
  XOR2_X1 U69 ( .A(n248), .B(n252), .Z(n249) );
  INV_X4 U70 ( .A(n247), .ZN(n252) );
  NOR3_X1 U71 ( .A1(\U10/DATA1_1 ), .A2(\U10/DATA1_14 ), .A3(\U10/DATA1_15 ), 
        .ZN(n383) );
  NAND2_X1 U72 ( .A1(n264), .A2(n263), .ZN(n257) );
  INV_X1 U73 ( .A(n301), .ZN(n286) );
  NAND2_X2 U74 ( .A1(n285), .A2(n284), .ZN(n301) );
  NAND3_X1 U75 ( .A1(n277), .A2(n279), .A3(n278), .ZN(n266) );
  INV_X1 U76 ( .A(n357), .ZN(n358) );
  XNOR2_X1 U77 ( .A(\U10/DATA1_0 ), .B(\add_48/B[0] ), .ZN(n246) );
  XOR2_X1 U78 ( .A(n347), .B(n344), .Z(n345) );
  NOR3_X1 U79 ( .A1(n381), .A2(\U10/DATA1_19 ), .A3(\U10/DATA1_0 ), .ZN(n382)
         );
  NAND2_X1 U80 ( .A1(n312), .A2(n311), .ZN(n306) );
  XOR2_X1 U81 ( .A(n330), .B(n326), .Z(n327) );
  XOR2_X1 U82 ( .A(n324), .B(n320), .Z(n321) );
  XOR2_X1 U83 ( .A(n342), .B(n338), .Z(n339) );
  XOR2_X1 U84 ( .A(n354), .B(n350), .Z(n351) );
  OAI21_X2 U85 ( .B1(n354), .B2(n353), .A(n352), .ZN(n357) );
  NAND2_X2 U86 ( .A1(StartIn), .A2(n239), .ZN(n240) );
  NAND2_X2 U87 ( .A1(StartIn), .A2(n238), .ZN(n241) );
  NOR2_X2 U88 ( .A1(n246), .A2(n362), .ZN(\U4/Z_0 ) );
  OAI22_X2 U89 ( .A1(n41), .A2(n238), .B1(n21), .B2(n240), .ZN(n81) );
  XOR2_X2 U90 ( .A(n20), .B(\add_48/B[1] ), .Z(n248) );
  NAND2_X2 U91 ( .A1(\add_48/B[0] ), .A2(n237), .ZN(n247) );
  NOR2_X2 U92 ( .A1(n249), .A2(n362), .ZN(\U4/Z_1 ) );
  OAI22_X2 U93 ( .A1(n40), .A2(n239), .B1(n20), .B2(n241), .ZN(n80) );
  INV_X4 U94 ( .A(\add_48/B[1] ), .ZN(n250) );
  NAND2_X2 U95 ( .A1(n20), .A2(n250), .ZN(n251) );
  NOR2_X2 U96 ( .A1(n254), .A2(n362), .ZN(\U4/Z_2 ) );
  OAI22_X2 U97 ( .A1(n39), .A2(n43), .B1(n256), .B2(n44), .ZN(n79) );
  NAND2_X2 U98 ( .A1(\add_48/B[2] ), .A2(\U10/DATA1_2 ), .ZN(n265) );
  INV_X4 U99 ( .A(\add_48/B[2] ), .ZN(n255) );
  NAND2_X2 U100 ( .A1(n256), .A2(n255), .ZN(n278) );
  NAND2_X2 U101 ( .A1(n278), .A2(n257), .ZN(n258) );
  NAND2_X2 U102 ( .A1(n265), .A2(n258), .ZN(n259) );
  NOR2_X2 U103 ( .A1(n260), .A2(n362), .ZN(\U4/Z_3 ) );
  OAI22_X2 U104 ( .A1(n38), .A2(n238), .B1(n262), .B2(n240), .ZN(n78) );
  INV_X4 U105 ( .A(\add_48/B[3] ), .ZN(n261) );
  NAND2_X2 U106 ( .A1(n262), .A2(n261), .ZN(n277) );
  NAND3_X2 U107 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n279) );
  NAND2_X2 U108 ( .A1(\add_48/B[3] ), .A2(\U10/DATA1_3 ), .ZN(n280) );
  NAND2_X2 U109 ( .A1(n266), .A2(n280), .ZN(n270) );
  NOR2_X2 U110 ( .A1(n268), .A2(n362), .ZN(\U4/Z_4 ) );
  OAI22_X2 U111 ( .A1(n37), .A2(n239), .B1(n17), .B2(n241), .ZN(n77) );
  XOR2_X2 U112 ( .A(\add_48/B[5] ), .B(\U10/DATA1_5 ), .Z(n273) );
  INV_X4 U113 ( .A(\add_48/B[4] ), .ZN(n269) );
  NAND2_X2 U114 ( .A1(n17), .A2(n269), .ZN(n275) );
  NAND2_X2 U115 ( .A1(n275), .A2(n270), .ZN(n271) );
  NAND2_X2 U116 ( .A1(n281), .A2(n271), .ZN(n272) );
  XNOR2_X2 U117 ( .A(n273), .B(n272), .ZN(n274) );
  NOR2_X2 U118 ( .A1(n274), .A2(n362), .ZN(\U4/Z_5 ) );
  OAI22_X2 U119 ( .A1(n36), .A2(n43), .B1(n16), .B2(n44), .ZN(n76) );
  INV_X4 U120 ( .A(n276), .ZN(n283) );
  NAND4_X2 U121 ( .A1(n283), .A2(n279), .A3(n278), .A4(n277), .ZN(n285) );
  NAND2_X2 U122 ( .A1(n281), .A2(n280), .ZN(n282) );
  NAND2_X2 U123 ( .A1(n283), .A2(n282), .ZN(n284) );
  NAND2_X2 U124 ( .A1(\add_48/B[5] ), .A2(\U10/DATA1_5 ), .ZN(n295) );
  NAND2_X2 U125 ( .A1(n286), .A2(n295), .ZN(n291) );
  NOR2_X2 U126 ( .A1(n288), .A2(n362), .ZN(\U4/Z_6 ) );
  OAI22_X2 U127 ( .A1(n35), .A2(n238), .B1(n290), .B2(n240), .ZN(n75) );
  NAND2_X2 U128 ( .A1(\add_48/B[6] ), .A2(\U10/DATA1_6 ), .ZN(n296) );
  INV_X4 U129 ( .A(\add_48/B[6] ), .ZN(n289) );
  NAND2_X2 U130 ( .A1(n290), .A2(n289), .ZN(n299) );
  NAND2_X2 U131 ( .A1(n299), .A2(n291), .ZN(n292) );
  NAND2_X2 U132 ( .A1(n296), .A2(n292), .ZN(n293) );
  NOR2_X2 U133 ( .A1(n294), .A2(n362), .ZN(\U4/Z_7 ) );
  OAI22_X2 U134 ( .A1(n34), .A2(n239), .B1(n298), .B2(n241), .ZN(n74) );
  NAND2_X2 U135 ( .A1(\add_48/B[7] ), .A2(\U10/DATA1_7 ), .ZN(n312) );
  NAND2_X2 U136 ( .A1(n296), .A2(n295), .ZN(n302) );
  INV_X4 U137 ( .A(\add_48/B[7] ), .ZN(n297) );
  NAND2_X2 U138 ( .A1(n298), .A2(n297), .ZN(n300) );
  NOR2_X2 U139 ( .A1(n304), .A2(n362), .ZN(\U4/Z_8 ) );
  OAI22_X2 U140 ( .A1(n33), .A2(n43), .B1(n385), .B2(n44), .ZN(n73) );
  XOR2_X2 U141 ( .A(\add_48/B[9] ), .B(\U10/DATA1_9 ), .Z(n309) );
  NAND2_X2 U142 ( .A1(\add_48/B[8] ), .A2(\U10/DATA1_8 ), .ZN(n313) );
  INV_X4 U143 ( .A(\add_48/B[8] ), .ZN(n305) );
  NAND2_X2 U144 ( .A1(n385), .A2(n305), .ZN(n314) );
  NAND2_X2 U145 ( .A1(n314), .A2(n306), .ZN(n307) );
  NAND2_X2 U146 ( .A1(n313), .A2(n307), .ZN(n308) );
  XNOR2_X2 U147 ( .A(n309), .B(n308), .ZN(n310) );
  NOR2_X2 U148 ( .A1(n310), .A2(n362), .ZN(\U4/Z_9 ) );
  OAI22_X2 U149 ( .A1(n32), .A2(n238), .B1(n384), .B2(n240), .ZN(n72) );
  NAND2_X2 U150 ( .A1(\add_48/B[9] ), .A2(\U10/DATA1_9 ), .ZN(n316) );
  NAND2_X2 U151 ( .A1(n316), .A2(n315), .ZN(n319) );
  XOR2_X2 U152 ( .A(\add_48/B[10] ), .B(\U10/DATA1_10 ), .Z(n317) );
  XOR2_X2 U153 ( .A(n221), .B(n317), .Z(n318) );
  NOR2_X2 U154 ( .A1(n318), .A2(n362), .ZN(\U4/Z_10 ) );
  OAI22_X2 U155 ( .A1(n31), .A2(n239), .B1(n11), .B2(n241), .ZN(n71) );
  XOR2_X2 U156 ( .A(\add_48/B[11] ), .B(\U10/DATA1_11 ), .Z(n320) );
  NOR2_X2 U157 ( .A1(n321), .A2(n362), .ZN(\U4/Z_11 ) );
  OAI22_X2 U158 ( .A1(n30), .A2(n43), .B1(n323), .B2(n44), .ZN(n70) );
  INV_X4 U159 ( .A(\add_48/B[11] ), .ZN(n322) );
  NAND2_X2 U160 ( .A1(n323), .A2(n322), .ZN(n325) );
  AOI22_X4 U161 ( .A1(n220), .A2(n325), .B1(\U10/DATA1_11 ), .B2(
        \add_48/B[11] ), .ZN(n330) );
  XOR2_X2 U162 ( .A(\add_48/B[12] ), .B(\U10/DATA1_12 ), .Z(n326) );
  NOR2_X2 U163 ( .A1(n327), .A2(n362), .ZN(\U4/Z_12 ) );
  OAI22_X2 U164 ( .A1(n29), .A2(n238), .B1(n329), .B2(n240), .ZN(n69) );
  INV_X4 U165 ( .A(\add_48/B[12] ), .ZN(n328) );
  NAND2_X2 U166 ( .A1(n329), .A2(n328), .ZN(n332) );
  INV_X4 U167 ( .A(n330), .ZN(n331) );
  XOR2_X2 U168 ( .A(\add_48/B[13] ), .B(\U10/DATA1_13 ), .Z(n333) );
  NOR2_X2 U169 ( .A1(n334), .A2(n362), .ZN(\U4/Z_13 ) );
  OAI22_X2 U170 ( .A1(n28), .A2(n239), .B1(n336), .B2(n241), .ZN(n68) );
  INV_X4 U171 ( .A(\add_48/B[13] ), .ZN(n335) );
  XOR2_X2 U172 ( .A(\add_48/B[14] ), .B(\U10/DATA1_14 ), .Z(n338) );
  NOR2_X2 U173 ( .A1(n339), .A2(n362), .ZN(\U4/Z_14 ) );
  OAI22_X2 U174 ( .A1(n27), .A2(n43), .B1(n341), .B2(n44), .ZN(n67) );
  INV_X4 U175 ( .A(\add_48/B[14] ), .ZN(n340) );
  NAND2_X2 U176 ( .A1(n341), .A2(n340), .ZN(n343) );
  AOI22_X4 U177 ( .A1(n224), .A2(n343), .B1(\U10/DATA1_14 ), .B2(
        \add_48/B[14] ), .ZN(n347) );
  XOR2_X2 U178 ( .A(\add_48/B[15] ), .B(\U10/DATA1_15 ), .Z(n344) );
  NOR2_X2 U179 ( .A1(n345), .A2(n362), .ZN(\U4/Z_15 ) );
  OAI22_X2 U180 ( .A1(n26), .A2(n238), .B1(n6), .B2(n240), .ZN(n66) );
  INV_X4 U181 ( .A(\add_48/B[15] ), .ZN(n346) );
  NAND2_X2 U182 ( .A1(n6), .A2(n346), .ZN(n349) );
  INV_X4 U183 ( .A(n347), .ZN(n348) );
  XOR2_X2 U184 ( .A(\add_48/B[16] ), .B(\U10/DATA1_16 ), .Z(n350) );
  NOR2_X2 U185 ( .A1(n351), .A2(n362), .ZN(\U4/Z_16 ) );
  OAI22_X2 U186 ( .A1(n25), .A2(n239), .B1(n5), .B2(n241), .ZN(n65) );
  NOR2_X2 U187 ( .A1(\add_48/B[16] ), .A2(\U10/DATA1_16 ), .ZN(n353) );
  NAND2_X2 U188 ( .A1(\add_48/B[16] ), .A2(\U10/DATA1_16 ), .ZN(n352) );
  NOR2_X2 U189 ( .A1(n355), .A2(n362), .ZN(\U4/Z_17 ) );
  OAI22_X2 U190 ( .A1(n24), .A2(n43), .B1(n380), .B2(n44), .ZN(n64) );
  XOR2_X2 U191 ( .A(n379), .B(\add_48/B[18] ), .Z(n361) );
  INV_X4 U192 ( .A(\add_48/B[17] ), .ZN(n356) );
  NAND2_X2 U193 ( .A1(n380), .A2(n356), .ZN(n359) );
  NAND2_X2 U194 ( .A1(n359), .A2(n357), .ZN(n368) );
  NAND2_X2 U195 ( .A1(\add_48/B[17] ), .A2(\U10/DATA1_17 ), .ZN(n369) );
  NOR2_X2 U196 ( .A1(n361), .A2(n369), .ZN(n363) );
  OAI22_X2 U197 ( .A1(n23), .A2(n238), .B1(n379), .B2(n240), .ZN(n63) );
  INV_X4 U198 ( .A(\add_48/B[18] ), .ZN(n365) );
  NAND2_X2 U199 ( .A1(n379), .A2(n365), .ZN(n372) );
  INV_X4 U200 ( .A(n372), .ZN(n367) );
  XOR2_X2 U201 ( .A(n366), .B(\add_48/B[19] ), .Z(n371) );
  NOR2_X2 U202 ( .A1(n367), .A2(n371), .ZN(n378) );
  NAND2_X2 U203 ( .A1(n369), .A2(n368), .ZN(n377) );
  NAND2_X2 U204 ( .A1(\add_48/B[18] ), .A2(\U10/DATA1_18 ), .ZN(n370) );
  NAND2_X2 U205 ( .A1(n371), .A2(n370), .ZN(n373) );
  OAI22_X2 U206 ( .A1(n22), .A2(n239), .B1(n366), .B2(n241), .ZN(n62) );
  NAND3_X2 U207 ( .A1(n5), .A2(n380), .A3(n379), .ZN(n381) );
  NAND4_X2 U208 ( .A1(n385), .A2(n384), .A3(n383), .A4(n382), .ZN(n390) );
  NOR3_X2 U209 ( .A1(\U10/DATA1_4 ), .A2(\U10/DATA1_2 ), .A3(\U10/DATA1_3 ), 
        .ZN(n388) );
  NAND3_X2 U210 ( .A1(n11), .A2(n298), .A3(n323), .ZN(n386) );
  NOR3_X2 U211 ( .A1(n386), .A2(\U10/DATA1_12 ), .A3(\U10/DATA1_13 ), .ZN(n387) );
  NAND4_X2 U212 ( .A1(n290), .A2(n16), .A3(n388), .A4(n387), .ZN(n389) );
  NOR2_X2 U213 ( .A1(n390), .A2(n389), .ZN(n391) );
  NOR3_X2 U214 ( .A1(n45), .A2(n362), .A3(n391), .ZN(\U8/Z_0 ) );
endmodule


module Cdf_Store ( clock, reset_n, StartIn, ResultIn, StoreAddressIn, WriteBus, 
        WriteAddress, WriteEnable );
  input [19:0] ResultIn;
  input [15:0] StoreAddressIn;
  output [127:0] WriteBus;
  output [15:0] WriteAddress;
  input clock, reset_n, StartIn;
  output WriteEnable;
  wire   n58, n57, n56, n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, n45,
         n44, n43, n42, n41, n40, n39, n182, n181, n180, n179, n178, n177,
         n176, n175, n174, n173, n172, n171, n170, n169, n168, n167, \U5/Z_0 ,
         \U5/Z_1 , \U5/Z_2 , \U5/Z_3 , \U5/Z_4 , \U5/Z_5 , \U5/Z_6 , \U5/Z_7 ,
         \U5/Z_8 , \U5/Z_9 , \U5/Z_10 , \U5/Z_11 , \U5/Z_12 , \U5/Z_13 ,
         \U5/Z_14 , \U5/Z_15 , \U5/Z_16 , \U5/Z_17 , \U5/Z_18 , \U5/Z_19 ,
         \U5/DATA1_0 , \U5/DATA1_1 , \U5/DATA1_2 , \U5/DATA1_3 , \U5/DATA1_4 ,
         \U5/DATA1_5 , \U5/DATA1_6 , \U5/DATA1_7 , \U5/DATA1_8 , \U5/DATA1_9 ,
         \U5/DATA1_10 , \U5/DATA1_11 , \U5/DATA1_12 , \U5/DATA1_13 ,
         \U5/DATA1_14 , \U5/DATA1_15 , \U5/DATA1_16 , \U5/DATA1_17 ,
         \U5/DATA1_18 , \U5/DATA1_19 , \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 ,
         \U4/Z_4 , \U4/Z_5 , \U4/Z_6 , \U4/Z_7 , \U4/Z_8 , \U4/Z_9 , \U4/Z_10 ,
         \U4/Z_11 , \U4/Z_12 , \U4/Z_13 , \U4/Z_14 , \U4/Z_15 , \U4/DATA1_0 ,
         \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 , \U4/DATA1_4 , \U4/DATA1_5 ,
         \U4/DATA1_6 , \U4/DATA1_7 , \U4/DATA1_8 , \U4/DATA1_9 , \U4/DATA1_10 ,
         \U4/DATA1_11 , \U4/DATA1_12 , \U4/DATA1_13 , \U4/DATA1_14 ,
         \U4/DATA1_15 , n517, n518, n519, n520, n521, n522, n523, n524, n525;
  assign \U5/DATA1_0  = ResultIn[0];
  assign \U5/DATA1_1  = ResultIn[1];
  assign \U5/DATA1_2  = ResultIn[2];
  assign \U5/DATA1_3  = ResultIn[3];
  assign \U5/DATA1_4  = ResultIn[4];
  assign \U5/DATA1_5  = ResultIn[5];
  assign \U5/DATA1_6  = ResultIn[6];
  assign \U5/DATA1_7  = ResultIn[7];
  assign \U5/DATA1_8  = ResultIn[8];
  assign \U5/DATA1_9  = ResultIn[9];
  assign \U5/DATA1_10  = ResultIn[10];
  assign \U5/DATA1_11  = ResultIn[11];
  assign \U5/DATA1_12  = ResultIn[12];
  assign \U5/DATA1_13  = ResultIn[13];
  assign \U5/DATA1_14  = ResultIn[14];
  assign \U5/DATA1_15  = ResultIn[15];
  assign \U5/DATA1_16  = ResultIn[16];
  assign \U5/DATA1_17  = ResultIn[17];
  assign \U5/DATA1_18  = ResultIn[18];
  assign \U5/DATA1_19  = ResultIn[19];
  assign \U4/DATA1_0  = StoreAddressIn[0];
  assign \U4/DATA1_1  = StoreAddressIn[1];
  assign \U4/DATA1_2  = StoreAddressIn[2];
  assign \U4/DATA1_3  = StoreAddressIn[3];
  assign \U4/DATA1_4  = StoreAddressIn[4];
  assign \U4/DATA1_5  = StoreAddressIn[5];
  assign \U4/DATA1_6  = StoreAddressIn[6];
  assign \U4/DATA1_7  = StoreAddressIn[7];
  assign \U4/DATA1_8  = StoreAddressIn[8];
  assign \U4/DATA1_9  = StoreAddressIn[9];
  assign \U4/DATA1_10  = StoreAddressIn[10];
  assign \U4/DATA1_11  = StoreAddressIn[11];
  assign \U4/DATA1_12  = StoreAddressIn[12];
  assign \U4/DATA1_13  = StoreAddressIn[13];
  assign \U4/DATA1_14  = StoreAddressIn[14];
  assign \U4/DATA1_15  = StoreAddressIn[15];

  TBUF_X2 \WriteBus_tri[0]  ( .A(n39), .EN(n525), .Z(WriteBus[0]) );
  TBUF_X2 \WriteBus_tri[1]  ( .A(n40), .EN(n519), .Z(WriteBus[1]) );
  TBUF_X2 \WriteBus_tri[2]  ( .A(n41), .EN(n519), .Z(WriteBus[2]) );
  TBUF_X2 \WriteBus_tri[3]  ( .A(n42), .EN(n519), .Z(WriteBus[3]) );
  TBUF_X2 \WriteBus_tri[4]  ( .A(n43), .EN(n520), .Z(WriteBus[4]) );
  TBUF_X2 \WriteBus_tri[5]  ( .A(n44), .EN(n520), .Z(WriteBus[5]) );
  TBUF_X2 \WriteBus_tri[6]  ( .A(n45), .EN(n520), .Z(WriteBus[6]) );
  TBUF_X2 \WriteBus_tri[7]  ( .A(n46), .EN(n525), .Z(WriteBus[7]) );
  TBUF_X2 \WriteBus_tri[8]  ( .A(n47), .EN(n518), .Z(WriteBus[8]) );
  TBUF_X2 \WriteBus_tri[9]  ( .A(n48), .EN(n518), .Z(WriteBus[9]) );
  TBUF_X2 \WriteBus_tri[10]  ( .A(n49), .EN(n518), .Z(WriteBus[10]) );
  TBUF_X2 \WriteBus_tri[11]  ( .A(n50), .EN(n518), .Z(WriteBus[11]) );
  TBUF_X2 \WriteBus_tri[12]  ( .A(n51), .EN(n520), .Z(WriteBus[12]) );
  TBUF_X2 \WriteBus_tri[13]  ( .A(n52), .EN(n519), .Z(WriteBus[13]) );
  TBUF_X2 \WriteBus_tri[14]  ( .A(n53), .EN(n525), .Z(WriteBus[14]) );
  TBUF_X2 \WriteBus_tri[15]  ( .A(n54), .EN(n519), .Z(WriteBus[15]) );
  TBUF_X2 \WriteBus_tri[16]  ( .A(n55), .EN(n519), .Z(WriteBus[16]) );
  TBUF_X2 \WriteBus_tri[17]  ( .A(n56), .EN(n519), .Z(WriteBus[17]) );
  TBUF_X2 \WriteBus_tri[18]  ( .A(n57), .EN(n518), .Z(WriteBus[18]) );
  TBUF_X2 \WriteBus_tri[19]  ( .A(n58), .EN(n519), .Z(WriteBus[19]) );
  TBUF_X2 \WriteBus_tri[20]  ( .A(1'b0), .EN(n519), .Z(WriteBus[20]) );
  TBUF_X2 \WriteBus_tri[21]  ( .A(1'b0), .EN(n525), .Z(WriteBus[21]) );
  TBUF_X2 \WriteBus_tri[22]  ( .A(1'b0), .EN(n519), .Z(WriteBus[22]) );
  TBUF_X2 \WriteBus_tri[23]  ( .A(1'b0), .EN(n520), .Z(WriteBus[23]) );
  TBUF_X2 \WriteBus_tri[24]  ( .A(1'b0), .EN(n519), .Z(WriteBus[24]) );
  TBUF_X2 \WriteBus_tri[25]  ( .A(1'b0), .EN(n520), .Z(WriteBus[25]) );
  TBUF_X2 \WriteBus_tri[26]  ( .A(1'b0), .EN(n519), .Z(WriteBus[26]) );
  TBUF_X2 \WriteBus_tri[27]  ( .A(1'b0), .EN(n518), .Z(WriteBus[27]) );
  TBUF_X2 \WriteBus_tri[28]  ( .A(1'b0), .EN(n519), .Z(WriteBus[28]) );
  TBUF_X2 \WriteBus_tri[29]  ( .A(1'b0), .EN(n525), .Z(WriteBus[29]) );
  TBUF_X2 \WriteBus_tri[30]  ( .A(1'b0), .EN(n519), .Z(WriteBus[30]) );
  TBUF_X2 \WriteBus_tri[31]  ( .A(1'b0), .EN(n519), .Z(WriteBus[31]) );
  TBUF_X2 \WriteBus_tri[32]  ( .A(1'b0), .EN(n520), .Z(WriteBus[32]) );
  TBUF_X2 \WriteBus_tri[33]  ( .A(1'b0), .EN(n519), .Z(WriteBus[33]) );
  TBUF_X2 \WriteBus_tri[34]  ( .A(1'b0), .EN(n520), .Z(WriteBus[34]) );
  TBUF_X2 \WriteBus_tri[35]  ( .A(1'b0), .EN(n519), .Z(WriteBus[35]) );
  TBUF_X2 \WriteBus_tri[36]  ( .A(1'b0), .EN(n520), .Z(WriteBus[36]) );
  TBUF_X2 \WriteBus_tri[37]  ( .A(1'b0), .EN(n525), .Z(WriteBus[37]) );
  TBUF_X2 \WriteBus_tri[38]  ( .A(1'b0), .EN(n518), .Z(WriteBus[38]) );
  TBUF_X2 \WriteBus_tri[39]  ( .A(1'b0), .EN(n519), .Z(WriteBus[39]) );
  TBUF_X2 \WriteBus_tri[40]  ( .A(1'b0), .EN(n518), .Z(WriteBus[40]) );
  TBUF_X2 \WriteBus_tri[41]  ( .A(1'b0), .EN(n520), .Z(WriteBus[41]) );
  TBUF_X2 \WriteBus_tri[42]  ( .A(1'b0), .EN(n519), .Z(WriteBus[42]) );
  TBUF_X2 \WriteBus_tri[43]  ( .A(1'b0), .EN(n518), .Z(WriteBus[43]) );
  TBUF_X2 \WriteBus_tri[44]  ( .A(1'b0), .EN(n519), .Z(WriteBus[44]) );
  TBUF_X2 \WriteBus_tri[45]  ( .A(1'b0), .EN(n519), .Z(WriteBus[45]) );
  TBUF_X2 \WriteBus_tri[46]  ( .A(1'b0), .EN(n525), .Z(WriteBus[46]) );
  TBUF_X2 \WriteBus_tri[47]  ( .A(1'b0), .EN(n520), .Z(WriteBus[47]) );
  TBUF_X2 \WriteBus_tri[48]  ( .A(1'b0), .EN(n518), .Z(WriteBus[48]) );
  TBUF_X2 \WriteBus_tri[49]  ( .A(1'b0), .EN(n518), .Z(WriteBus[49]) );
  TBUF_X2 \WriteBus_tri[50]  ( .A(1'b0), .EN(n519), .Z(WriteBus[50]) );
  TBUF_X2 \WriteBus_tri[51]  ( .A(1'b0), .EN(n518), .Z(WriteBus[51]) );
  TBUF_X2 \WriteBus_tri[52]  ( .A(1'b0), .EN(n520), .Z(WriteBus[52]) );
  TBUF_X2 \WriteBus_tri[53]  ( .A(1'b0), .EN(n518), .Z(WriteBus[53]) );
  TBUF_X2 \WriteBus_tri[54]  ( .A(1'b0), .EN(n518), .Z(WriteBus[54]) );
  TBUF_X2 \WriteBus_tri[55]  ( .A(1'b0), .EN(n519), .Z(WriteBus[55]) );
  TBUF_X2 \WriteBus_tri[56]  ( .A(1'b0), .EN(n519), .Z(WriteBus[56]) );
  TBUF_X2 \WriteBus_tri[57]  ( .A(1'b0), .EN(n520), .Z(WriteBus[57]) );
  TBUF_X2 \WriteBus_tri[58]  ( .A(1'b0), .EN(n519), .Z(WriteBus[58]) );
  TBUF_X2 \WriteBus_tri[59]  ( .A(1'b0), .EN(n520), .Z(WriteBus[59]) );
  TBUF_X2 \WriteBus_tri[60]  ( .A(1'b0), .EN(n520), .Z(WriteBus[60]) );
  TBUF_X2 \WriteBus_tri[61]  ( .A(1'b0), .EN(n518), .Z(WriteBus[61]) );
  TBUF_X2 \WriteBus_tri[62]  ( .A(1'b0), .EN(n520), .Z(WriteBus[62]) );
  TBUF_X2 \WriteBus_tri[63]  ( .A(1'b0), .EN(n520), .Z(WriteBus[63]) );
  TBUF_X2 \WriteBus_tri[64]  ( .A(1'b0), .EN(n520), .Z(WriteBus[64]) );
  TBUF_X2 \WriteBus_tri[65]  ( .A(1'b0), .EN(n519), .Z(WriteBus[65]) );
  TBUF_X2 \WriteBus_tri[66]  ( .A(1'b0), .EN(n520), .Z(WriteBus[66]) );
  TBUF_X2 \WriteBus_tri[67]  ( .A(1'b0), .EN(n520), .Z(WriteBus[67]) );
  TBUF_X2 \WriteBus_tri[68]  ( .A(1'b0), .EN(n520), .Z(WriteBus[68]) );
  TBUF_X2 \WriteBus_tri[69]  ( .A(1'b0), .EN(n520), .Z(WriteBus[69]) );
  TBUF_X2 \WriteBus_tri[70]  ( .A(1'b0), .EN(n520), .Z(WriteBus[70]) );
  TBUF_X2 \WriteBus_tri[71]  ( .A(1'b0), .EN(n520), .Z(WriteBus[71]) );
  TBUF_X2 \WriteBus_tri[72]  ( .A(1'b0), .EN(n518), .Z(WriteBus[72]) );
  TBUF_X2 \WriteBus_tri[73]  ( .A(1'b0), .EN(n520), .Z(WriteBus[73]) );
  TBUF_X2 \WriteBus_tri[74]  ( .A(1'b0), .EN(n525), .Z(WriteBus[74]) );
  TBUF_X2 \WriteBus_tri[75]  ( .A(1'b0), .EN(n520), .Z(WriteBus[75]) );
  TBUF_X2 \WriteBus_tri[76]  ( .A(1'b0), .EN(n519), .Z(WriteBus[76]) );
  TBUF_X2 \WriteBus_tri[77]  ( .A(1'b0), .EN(n520), .Z(WriteBus[77]) );
  TBUF_X2 \WriteBus_tri[78]  ( .A(1'b0), .EN(n520), .Z(WriteBus[78]) );
  TBUF_X2 \WriteBus_tri[79]  ( .A(1'b0), .EN(n525), .Z(WriteBus[79]) );
  TBUF_X2 \WriteBus_tri[80]  ( .A(1'b0), .EN(n518), .Z(WriteBus[80]) );
  TBUF_X2 \WriteBus_tri[81]  ( .A(1'b0), .EN(n519), .Z(WriteBus[81]) );
  TBUF_X2 \WriteBus_tri[82]  ( .A(1'b0), .EN(n520), .Z(WriteBus[82]) );
  TBUF_X2 \WriteBus_tri[83]  ( .A(1'b0), .EN(n519), .Z(WriteBus[83]) );
  TBUF_X2 \WriteBus_tri[84]  ( .A(1'b0), .EN(n519), .Z(WriteBus[84]) );
  TBUF_X2 \WriteBus_tri[85]  ( .A(1'b0), .EN(n518), .Z(WriteBus[85]) );
  TBUF_X2 \WriteBus_tri[86]  ( .A(1'b0), .EN(n518), .Z(WriteBus[86]) );
  TBUF_X2 \WriteBus_tri[87]  ( .A(1'b0), .EN(n520), .Z(WriteBus[87]) );
  TBUF_X2 \WriteBus_tri[88]  ( .A(1'b0), .EN(n518), .Z(WriteBus[88]) );
  TBUF_X2 \WriteBus_tri[89]  ( .A(1'b0), .EN(n520), .Z(WriteBus[89]) );
  TBUF_X2 \WriteBus_tri[90]  ( .A(1'b0), .EN(n518), .Z(WriteBus[90]) );
  TBUF_X2 \WriteBus_tri[91]  ( .A(1'b0), .EN(n518), .Z(WriteBus[91]) );
  TBUF_X2 \WriteBus_tri[92]  ( .A(1'b0), .EN(n525), .Z(WriteBus[92]) );
  TBUF_X2 \WriteBus_tri[93]  ( .A(1'b0), .EN(n520), .Z(WriteBus[93]) );
  TBUF_X2 \WriteBus_tri[94]  ( .A(1'b0), .EN(n519), .Z(WriteBus[94]) );
  TBUF_X2 \WriteBus_tri[95]  ( .A(1'b0), .EN(n518), .Z(WriteBus[95]) );
  TBUF_X2 \WriteBus_tri[96]  ( .A(1'b0), .EN(n520), .Z(WriteBus[96]) );
  TBUF_X2 \WriteBus_tri[97]  ( .A(1'b0), .EN(n519), .Z(WriteBus[97]) );
  TBUF_X2 \WriteBus_tri[98]  ( .A(1'b0), .EN(n519), .Z(WriteBus[98]) );
  TBUF_X2 \WriteBus_tri[99]  ( .A(1'b0), .EN(n518), .Z(WriteBus[99]) );
  TBUF_X2 \WriteBus_tri[100]  ( .A(1'b0), .EN(n520), .Z(WriteBus[100]) );
  TBUF_X2 \WriteBus_tri[101]  ( .A(1'b0), .EN(n525), .Z(WriteBus[101]) );
  TBUF_X2 \WriteBus_tri[102]  ( .A(1'b0), .EN(n518), .Z(WriteBus[102]) );
  TBUF_X2 \WriteBus_tri[103]  ( .A(1'b0), .EN(n525), .Z(WriteBus[103]) );
  TBUF_X2 \WriteBus_tri[104]  ( .A(1'b0), .EN(n525), .Z(WriteBus[104]) );
  TBUF_X2 \WriteBus_tri[105]  ( .A(1'b0), .EN(n525), .Z(WriteBus[105]) );
  TBUF_X2 \WriteBus_tri[106]  ( .A(1'b0), .EN(n519), .Z(WriteBus[106]) );
  TBUF_X2 \WriteBus_tri[107]  ( .A(1'b0), .EN(n518), .Z(WriteBus[107]) );
  TBUF_X2 \WriteBus_tri[108]  ( .A(1'b0), .EN(n520), .Z(WriteBus[108]) );
  TBUF_X2 \WriteBus_tri[109]  ( .A(1'b0), .EN(n518), .Z(WriteBus[109]) );
  TBUF_X2 \WriteBus_tri[110]  ( .A(1'b0), .EN(n518), .Z(WriteBus[110]) );
  TBUF_X2 \WriteBus_tri[111]  ( .A(1'b0), .EN(n525), .Z(WriteBus[111]) );
  TBUF_X2 \WriteBus_tri[112]  ( .A(1'b0), .EN(n518), .Z(WriteBus[112]) );
  TBUF_X2 \WriteBus_tri[113]  ( .A(1'b0), .EN(n519), .Z(WriteBus[113]) );
  TBUF_X2 \WriteBus_tri[114]  ( .A(1'b0), .EN(n518), .Z(WriteBus[114]) );
  TBUF_X2 \WriteBus_tri[115]  ( .A(1'b0), .EN(n519), .Z(WriteBus[115]) );
  TBUF_X2 \WriteBus_tri[116]  ( .A(1'b0), .EN(n518), .Z(WriteBus[116]) );
  TBUF_X2 \WriteBus_tri[117]  ( .A(1'b0), .EN(n520), .Z(WriteBus[117]) );
  TBUF_X2 \WriteBus_tri[118]  ( .A(1'b0), .EN(n518), .Z(WriteBus[118]) );
  TBUF_X2 \WriteBus_tri[119]  ( .A(1'b0), .EN(n520), .Z(WriteBus[119]) );
  TBUF_X2 \WriteBus_tri[120]  ( .A(1'b0), .EN(n518), .Z(WriteBus[120]) );
  TBUF_X2 \WriteBus_tri[121]  ( .A(1'b0), .EN(n518), .Z(WriteBus[121]) );
  TBUF_X2 \WriteBus_tri[122]  ( .A(1'b0), .EN(n525), .Z(WriteBus[122]) );
  TBUF_X2 \WriteBus_tri[123]  ( .A(1'b0), .EN(n518), .Z(WriteBus[123]) );
  TBUF_X2 \WriteBus_tri[124]  ( .A(1'b0), .EN(n519), .Z(WriteBus[124]) );
  TBUF_X2 \WriteBus_tri[125]  ( .A(1'b0), .EN(n518), .Z(WriteBus[125]) );
  TBUF_X2 \WriteBus_tri[126]  ( .A(1'b0), .EN(n518), .Z(WriteBus[126]) );
  TBUF_X2 \WriteBus_tri[127]  ( .A(1'b0), .EN(n518), .Z(WriteBus[127]) );
  TBUF_X2 \WriteAddress_tri[0]  ( .A(n167), .EN(n525), .Z(WriteAddress[0]) );
  TBUF_X2 \WriteAddress_tri[1]  ( .A(n168), .EN(n520), .Z(WriteAddress[1]) );
  TBUF_X2 \WriteAddress_tri[2]  ( .A(n169), .EN(n525), .Z(WriteAddress[2]) );
  TBUF_X2 \WriteAddress_tri[3]  ( .A(n170), .EN(n518), .Z(WriteAddress[3]) );
  TBUF_X2 \WriteAddress_tri[4]  ( .A(n171), .EN(n525), .Z(WriteAddress[4]) );
  TBUF_X2 \WriteAddress_tri[5]  ( .A(n172), .EN(n525), .Z(WriteAddress[5]) );
  TBUF_X2 \WriteAddress_tri[6]  ( .A(n173), .EN(n525), .Z(WriteAddress[6]) );
  TBUF_X2 \WriteAddress_tri[7]  ( .A(n174), .EN(n519), .Z(WriteAddress[7]) );
  TBUF_X2 \WriteAddress_tri[8]  ( .A(n175), .EN(n525), .Z(WriteAddress[8]) );
  TBUF_X2 \WriteAddress_tri[9]  ( .A(n176), .EN(n518), .Z(WriteAddress[9]) );
  TBUF_X2 \WriteAddress_tri[10]  ( .A(n177), .EN(n525), .Z(WriteAddress[10])
         );
  TBUF_X2 \WriteAddress_tri[11]  ( .A(n178), .EN(n525), .Z(WriteAddress[11])
         );
  TBUF_X2 \WriteAddress_tri[12]  ( .A(n179), .EN(n519), .Z(WriteAddress[12])
         );
  TBUF_X2 \WriteAddress_tri[13]  ( .A(n180), .EN(n525), .Z(WriteAddress[13])
         );
  TBUF_X2 \WriteAddress_tri[14]  ( .A(n181), .EN(n520), .Z(WriteAddress[14])
         );
  TBUF_X2 \WriteAddress_tri[15]  ( .A(n182), .EN(n525), .Z(WriteAddress[15])
         );
  TBUF_X2 WriteEnable_tri ( .A(1'b1), .EN(n525), .Z(WriteEnable) );
  AND2_X1 U6 ( .A1(\U5/DATA1_9 ), .A2(StartIn), .ZN(\U5/Z_9 ) );
  AND2_X1 U7 ( .A1(\U5/DATA1_8 ), .A2(StartIn), .ZN(\U5/Z_8 ) );
  AND2_X1 U8 ( .A1(\U5/DATA1_7 ), .A2(StartIn), .ZN(\U5/Z_7 ) );
  AND2_X1 U9 ( .A1(\U5/DATA1_6 ), .A2(StartIn), .ZN(\U5/Z_6 ) );
  AND2_X1 U10 ( .A1(\U5/DATA1_5 ), .A2(StartIn), .ZN(\U5/Z_5 ) );
  AND2_X1 U12 ( .A1(\U5/DATA1_3 ), .A2(StartIn), .ZN(\U5/Z_3 ) );
  AND2_X1 U13 ( .A1(\U5/DATA1_2 ), .A2(StartIn), .ZN(\U5/Z_2 ) );
  AND2_X1 U14 ( .A1(\U5/DATA1_19 ), .A2(StartIn), .ZN(\U5/Z_19 ) );
  AND2_X1 U15 ( .A1(\U5/DATA1_18 ), .A2(StartIn), .ZN(\U5/Z_18 ) );
  AND2_X1 U16 ( .A1(\U5/DATA1_17 ), .A2(StartIn), .ZN(\U5/Z_17 ) );
  AND2_X1 U17 ( .A1(\U5/DATA1_16 ), .A2(StartIn), .ZN(\U5/Z_16 ) );
  AND2_X1 U18 ( .A1(\U5/DATA1_15 ), .A2(StartIn), .ZN(\U5/Z_15 ) );
  AND2_X1 U19 ( .A1(\U5/DATA1_14 ), .A2(StartIn), .ZN(\U5/Z_14 ) );
  AND2_X1 U20 ( .A1(\U5/DATA1_13 ), .A2(StartIn), .ZN(\U5/Z_13 ) );
  AND2_X1 U21 ( .A1(\U5/DATA1_12 ), .A2(StartIn), .ZN(\U5/Z_12 ) );
  AND2_X1 U22 ( .A1(\U5/DATA1_11 ), .A2(StartIn), .ZN(\U5/Z_11 ) );
  AND2_X1 U23 ( .A1(\U5/DATA1_10 ), .A2(StartIn), .ZN(\U5/Z_10 ) );
  AND2_X1 U24 ( .A1(\U5/DATA1_1 ), .A2(StartIn), .ZN(\U5/Z_1 ) );
  AND2_X1 U26 ( .A1(\U4/DATA1_9 ), .A2(StartIn), .ZN(\U4/Z_9 ) );
  AND2_X1 U27 ( .A1(\U4/DATA1_8 ), .A2(StartIn), .ZN(\U4/Z_8 ) );
  AND2_X1 U28 ( .A1(\U4/DATA1_7 ), .A2(StartIn), .ZN(\U4/Z_7 ) );
  AND2_X1 U29 ( .A1(\U4/DATA1_6 ), .A2(StartIn), .ZN(\U4/Z_6 ) );
  AND2_X1 U30 ( .A1(\U4/DATA1_5 ), .A2(StartIn), .ZN(\U4/Z_5 ) );
  AND2_X1 U31 ( .A1(\U4/DATA1_4 ), .A2(StartIn), .ZN(\U4/Z_4 ) );
  AND2_X1 U32 ( .A1(\U4/DATA1_3 ), .A2(StartIn), .ZN(\U4/Z_3 ) );
  AND2_X1 U33 ( .A1(\U4/DATA1_2 ), .A2(StartIn), .ZN(\U4/Z_2 ) );
  AND2_X1 U34 ( .A1(\U4/DATA1_15 ), .A2(StartIn), .ZN(\U4/Z_15 ) );
  AND2_X1 U35 ( .A1(\U4/DATA1_14 ), .A2(StartIn), .ZN(\U4/Z_14 ) );
  AND2_X1 U36 ( .A1(\U4/DATA1_13 ), .A2(StartIn), .ZN(\U4/Z_13 ) );
  AND2_X1 U37 ( .A1(\U4/DATA1_12 ), .A2(StartIn), .ZN(\U4/Z_12 ) );
  AND2_X1 U38 ( .A1(\U4/DATA1_11 ), .A2(StartIn), .ZN(\U4/Z_11 ) );
  AND2_X1 U39 ( .A1(\U4/DATA1_10 ), .A2(StartIn), .ZN(\U4/Z_10 ) );
  AND2_X1 U40 ( .A1(\U4/DATA1_1 ), .A2(StartIn), .ZN(\U4/Z_1 ) );
  AND2_X1 U41 ( .A1(\U4/DATA1_0 ), .A2(StartIn), .ZN(\U4/Z_0 ) );
  DFFR_X2 Write_reg ( .D(StartIn), .CK(clock), .RN(n522), .Q(n517), .QN(n525)
         );
  DFFR_X2 \Write_Bus_reg[19]  ( .D(\U5/Z_19 ), .CK(clock), .RN(reset_n), .Q(
        n58) );
  DFFR_X2 \Write_Bus_reg[18]  ( .D(\U5/Z_18 ), .CK(clock), .RN(n524), .Q(n57)
         );
  DFFR_X2 \Write_Bus_reg[17]  ( .D(\U5/Z_17 ), .CK(clock), .RN(n524), .Q(n56)
         );
  DFFR_X2 \Write_Bus_reg[16]  ( .D(\U5/Z_16 ), .CK(clock), .RN(n524), .Q(n55)
         );
  DFFR_X2 \Write_Bus_reg[15]  ( .D(\U5/Z_15 ), .CK(clock), .RN(n524), .Q(n54)
         );
  DFFR_X2 \Write_Bus_reg[14]  ( .D(\U5/Z_14 ), .CK(clock), .RN(n524), .Q(n53)
         );
  DFFR_X2 \Write_Bus_reg[13]  ( .D(\U5/Z_13 ), .CK(clock), .RN(n524), .Q(n52)
         );
  DFFR_X2 \Write_Bus_reg[12]  ( .D(\U5/Z_12 ), .CK(clock), .RN(n524), .Q(n51)
         );
  DFFR_X2 \Write_Bus_reg[11]  ( .D(\U5/Z_11 ), .CK(clock), .RN(n524), .Q(n50)
         );
  DFFR_X2 \Write_Bus_reg[10]  ( .D(\U5/Z_10 ), .CK(clock), .RN(n524), .Q(n49)
         );
  DFFR_X2 \Write_Bus_reg[9]  ( .D(\U5/Z_9 ), .CK(clock), .RN(n524), .Q(n48) );
  DFFR_X2 \Write_Bus_reg[8]  ( .D(\U5/Z_8 ), .CK(clock), .RN(n524), .Q(n47) );
  DFFR_X2 \Write_Bus_reg[7]  ( .D(\U5/Z_7 ), .CK(clock), .RN(n524), .Q(n46) );
  DFFR_X2 \Write_Bus_reg[6]  ( .D(\U5/Z_6 ), .CK(clock), .RN(n523), .Q(n45) );
  DFFR_X2 \Write_Bus_reg[5]  ( .D(\U5/Z_5 ), .CK(clock), .RN(n523), .Q(n44) );
  DFFR_X2 \Write_Bus_reg[3]  ( .D(\U5/Z_3 ), .CK(clock), .RN(n523), .Q(n42) );
  DFFR_X2 \Write_Bus_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .RN(n523), .Q(n41) );
  DFFR_X2 \Write_Bus_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .RN(n523), .Q(n40) );
  DFFR_X2 \WriteAddr_reg[15]  ( .D(\U4/Z_15 ), .CK(clock), .RN(n523), .Q(n182)
         );
  DFFR_X2 \WriteAddr_reg[14]  ( .D(\U4/Z_14 ), .CK(clock), .RN(n523), .Q(n181)
         );
  DFFR_X2 \WriteAddr_reg[13]  ( .D(\U4/Z_13 ), .CK(clock), .RN(n523), .Q(n180)
         );
  DFFR_X2 \WriteAddr_reg[12]  ( .D(\U4/Z_12 ), .CK(clock), .RN(n523), .Q(n179)
         );
  DFFR_X2 \WriteAddr_reg[11]  ( .D(\U4/Z_11 ), .CK(clock), .RN(n523), .Q(n178)
         );
  DFFR_X2 \WriteAddr_reg[10]  ( .D(\U4/Z_10 ), .CK(clock), .RN(n522), .Q(n177)
         );
  DFFR_X2 \WriteAddr_reg[9]  ( .D(\U4/Z_9 ), .CK(clock), .RN(n522), .Q(n176)
         );
  DFFR_X2 \WriteAddr_reg[8]  ( .D(\U4/Z_8 ), .CK(clock), .RN(n522), .Q(n175)
         );
  DFFR_X2 \WriteAddr_reg[7]  ( .D(\U4/Z_7 ), .CK(clock), .RN(n522), .Q(n174)
         );
  DFFR_X2 \WriteAddr_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n522), .Q(n173)
         );
  DFFR_X2 \WriteAddr_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n522), .Q(n172)
         );
  DFFR_X2 \WriteAddr_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(n522), .Q(n171)
         );
  DFFR_X2 \WriteAddr_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n522), .Q(n170)
         );
  DFFR_X2 \WriteAddr_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .RN(n522), .Q(n169)
         );
  DFFR_X2 \WriteAddr_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .RN(n522), .Q(n168)
         );
  DFFR_X2 \WriteAddr_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .RN(n522), .Q(n167)
         );
  DFFR_X2 \Write_Bus_reg[4]  ( .D(\U5/Z_4 ), .CK(clock), .RN(n523), .Q(n43) );
  DFFR_X2 \Write_Bus_reg[0]  ( .D(\U5/Z_0 ), .CK(clock), .RN(n523), .Q(n39) );
  INV_X4 U5 ( .A(n521), .ZN(n523) );
  INV_X4 U11 ( .A(n521), .ZN(n524) );
  INV_X4 U25 ( .A(n521), .ZN(n522) );
  INV_X4 U42 ( .A(reset_n), .ZN(n521) );
  INV_X4 U43 ( .A(n517), .ZN(n518) );
  INV_X4 U44 ( .A(n517), .ZN(n520) );
  INV_X4 U45 ( .A(n517), .ZN(n519) );
  AND2_X4 U46 ( .A1(\U5/DATA1_4 ), .A2(StartIn), .ZN(\U5/Z_4 ) );
  AND2_X4 U47 ( .A1(\U5/DATA1_0 ), .A2(StartIn), .ZN(\U5/Z_0 ) );
endmodule


module Cdf_top ( clock, reset_n, start, SP_ReadBus, SP_ReadAddress, 
        WriteEnable, Output_MEMBus, Output_MEMAddress, Cdf_Min, done, 
        input_base_offset, cdf_valid );
  input [127:0] SP_ReadBus;
  output [15:0] SP_ReadAddress;
  output [127:0] Output_MEMBus;
  output [15:0] Output_MEMAddress;
  output [19:0] Cdf_Min;
  input clock, reset_n, start, input_base_offset;
  output WriteEnable, done, cdf_valid;
  wire   start_to_accumlate, start_to_store, n1, n2;
  wire   [19:0] Accumlate;
  wire   [19:0] AccumlateResult;
  wire   [15:0] store_address;
  wire   [15:0] store_address_to_store;

  Cdf_Fetch stage1 ( .clock(clock), .reset_n(n1), .start(start), .ReadBus(
        SP_ReadBus), .ReadAddr(SP_ReadAddress), .AccumlateOut(Accumlate), 
        .StartOut(start_to_accumlate), .StoreAddress(store_address), 
        .input_base_offset(input_base_offset), .done(done) );
  Cdf_Accumlate stage2 ( .clock(clock), .reset_n(n1), .AccumlateIn(Accumlate), 
        .StartIn(start_to_accumlate), .StoreAddressIn(store_address), 
        .AccumlateResult(AccumlateResult), .StoreAddressOut(
        store_address_to_store), .StartOut(start_to_store), .CdfMin(Cdf_Min), 
        .CdfValid(cdf_valid) );
  Cdf_Store stage3 ( .clock(clock), .reset_n(n1), .StartIn(start_to_store), 
        .ResultIn(AccumlateResult), .StoreAddressIn(store_address_to_store), 
        .WriteBus(Output_MEMBus), .WriteAddress(Output_MEMAddress), 
        .WriteEnable(WriteEnable) );
  INV_X4 U1 ( .A(n2), .ZN(n1) );
  INV_X4 U2 ( .A(reset_n), .ZN(n2) );
endmodule


module input_pipeline ( start, clock, rst_n, m1ReadBus, m2ReadBus, 
        inputBaseOffset, m1ReadAddr, m2ReadAddr, m2WriteAddr, m3WriteAddr, 
        m2WriteBus, m3WriteBus, m2WE, m3WE, done, cdf_min, cdf_valid );
  input [127:0] m1ReadBus;
  input [127:0] m2ReadBus;
  output [15:0] m1ReadAddr;
  output [15:0] m2ReadAddr;
  output [15:0] m2WriteAddr;
  output [15:0] m3WriteAddr;
  output [127:0] m2WriteBus;
  output [127:0] m3WriteBus;
  output [19:0] cdf_min;
  input start, clock, rst_n, inputBaseOffset;
  output m2WE, m3WE, done, cdf_valid;
  wire   \U3/U1/Z_0 , \U3/U1/DATA2_35 , \U3/U1/DATA1_0 , \U3/U1/DATA1_1 ,
         \U3/U1/DATA1_2 , \U3/U1/DATA1_3 , \U3/U1/DATA1_4 , \U3/U1/DATA1_5 ,
         \U3/U1/DATA1_6 , \U3/U1/DATA1_7 , \U3/U1/DATA1_8 , \U3/U1/DATA1_9 ,
         \U3/U1/DATA1_10 , \U3/U1/DATA1_11 , \U3/U1/DATA1_12 ,
         \U3/U1/DATA1_13 , \U3/U1/DATA1_14 , \U3/U1/DATA1_15 ,
         \U3/U1/DATA1_16 , \U3/U1/DATA1_17 , \U3/U1/DATA1_18 ,
         \U3/U1/DATA1_19 , \U3/U1/DATA1_20 , \U3/U1/DATA1_21 ,
         \U3/U1/DATA1_22 , \U3/U1/DATA1_23 , \U3/U1/DATA1_24 ,
         \U3/U1/DATA1_25 , \U3/U1/DATA1_26 , \U3/U1/DATA1_27 ,
         \U3/U1/DATA1_28 , \U3/U1/DATA1_29 , \U3/U1/DATA1_30 ,
         \U3/U1/DATA1_31 , \U3/U1/DATA1_32 , \U3/U1/DATA1_33 ,
         \U3/U1/DATA1_34 , \U3/U1/DATA1_35 , \U36/DATA2_0 , \U36/DATA2_1 ,
         \U36/DATA2_2 , \U36/DATA2_3 , \U36/DATA2_4 , \U36/DATA2_5 ,
         \U36/DATA2_6 , \U36/DATA2_7 , \U36/DATA2_8 , \U36/DATA2_9 ,
         \U36/DATA2_10 , \U36/DATA2_11 , \U36/DATA2_12 , \U36/DATA2_13 ,
         \U36/DATA2_14 , \U36/DATA2_15 , \U36/DATA2_16 , \U36/DATA2_17 ,
         \U36/DATA2_18 , \U36/DATA2_19 , \U36/DATA2_20 , \U36/DATA2_21 ,
         \U36/DATA2_22 , \U36/DATA2_23 , \U36/DATA2_24 , \U36/DATA2_25 ,
         \U36/DATA2_26 , \U36/DATA2_27 , \U36/DATA2_28 , \U36/DATA2_29 ,
         \U36/DATA2_30 , \U36/DATA2_31 , \U36/DATA2_32 , \U36/DATA2_33 ,
         \U36/DATA2_34 , \U36/DATA2_35 , \U36/DATA2_36 , \U36/DATA2_37 ,
         \U36/DATA2_38 , \U36/DATA2_39 , \U36/DATA2_40 , \U36/DATA2_41 ,
         \U36/DATA2_42 , \U36/DATA2_43 , \U36/DATA2_44 , \U36/DATA2_45 ,
         \U36/DATA2_46 , \U36/DATA2_47 , \U36/DATA2_48 , \U36/DATA2_49 ,
         \U36/DATA2_50 , \U36/DATA2_51 , \U36/DATA2_52 , \U36/DATA2_53 ,
         \U36/DATA2_54 , \U36/DATA2_55 , \U36/DATA2_56 , \U36/DATA2_57 ,
         \U36/DATA2_58 , \U36/DATA2_59 , \U36/DATA2_60 , \U36/DATA2_61 ,
         \U36/DATA2_62 , \U36/DATA2_63 , \U36/DATA2_64 , \U36/DATA2_65 ,
         \U36/DATA2_66 , \U36/DATA2_67 , \U36/DATA2_68 , \U36/DATA2_69 ,
         \U36/DATA2_70 , \U36/DATA1_7 , \U36/DATA1_8 , \U36/DATA1_9 ,
         \U36/DATA1_10 , \U36/DATA1_11 , \U36/DATA1_12 , \U36/DATA1_13 ,
         \U36/DATA1_14 , \U36/DATA1_15 , \U36/DATA1_16 , \U36/DATA1_17 ,
         \U36/DATA1_18 , \U36/DATA1_19 , \U36/DATA1_20 , \U36/DATA1_21 ,
         \U36/DATA1_22 , \U36/DATA1_23 , \U36/DATA1_24 , \U36/DATA1_25 ,
         \U36/DATA1_26 , \U36/DATA1_27 , \U36/DATA1_28 , \U36/DATA1_29 ,
         \U36/DATA1_30 , \U36/DATA1_31 , \U36/DATA1_32 , \U36/DATA1_33 ,
         \U36/DATA1_34 , \U36/DATA1_35 , \U36/DATA1_36 , \U36/DATA1_37 ,
         \U36/DATA1_38 , \U36/DATA1_39 , \U36/DATA1_40 , \U36/DATA1_41 ,
         \U36/DATA1_42 , \U36/DATA1_43 , \U36/DATA1_44 , \U36/DATA1_45 ,
         \U36/DATA1_46 , \U36/DATA1_47 , \U36/DATA1_48 , \U36/DATA1_49 ,
         \U36/DATA1_50 , \U36/DATA1_51 , \U36/DATA1_52 , \U36/DATA1_53 ,
         \U36/DATA1_54 , \U36/DATA1_55 , \U36/DATA1_56 , \U36/DATA1_57 ,
         \U36/DATA1_58 , \U36/DATA1_59 , \U36/DATA1_60 , \U36/DATA1_61 ,
         \U36/DATA1_62 , \U36/DATA1_63 , \U29/Z_0 , \U29/Z_1 , \U29/Z_2 ,
         \U29/Z_3 , \U29/Z_4 , \U29/Z_5 , \U29/Z_6 , \U29/Z_7 , \U29/DATA2_0 ,
         \U29/DATA2_1 , \U29/DATA1_0 , \U29/DATA1_1 , \U29/DATA1_2 ,
         \U29/DATA1_3 , \U29/DATA1_4 , \U29/DATA1_5 , \U29/DATA1_6 ,
         \U29/DATA1_7 , \U29/DATA1_8 , \U29/DATA1_9 , \U29/DATA1_10 ,
         \U29/DATA1_11 , \U29/DATA1_12 , \U29/DATA1_13 , \U29/DATA1_14 ,
         \U29/DATA1_15 , \U28/Z_0 , \U28/DATA1_0 , \U27/Z_0 , \U27/Z_1 ,
         \U27/Z_2 , \U27/Z_3 , \U27/Z_4 , \U27/Z_5 , \U27/Z_6 , \U27/Z_7 ,
         \U27/DATA2_0 , \U27/DATA2_1 , \U27/DATA2_2 , \U27/DATA2_3 ,
         \U27/DATA2_4 , \U27/DATA2_5 , \U27/DATA2_6 , \U27/DATA2_7 ,
         \U27/DATA1_0 , \U27/DATA1_1 , \U27/DATA1_2 , \U27/DATA1_3 ,
         \U27/DATA1_4 , \U27/DATA1_5 , \U27/DATA1_6 , \U27/DATA1_7 ,
         \U27/DATA1_8 , \U27/DATA1_9 , \U27/DATA1_10 , \U27/DATA1_11 ,
         \U27/DATA1_12 , \U27/DATA1_13 , \U27/DATA1_14 , \U27/DATA1_15 ,
         \U26/Z_0 , \U26/Z_1 , \U26/Z_2 , \U26/Z_3 , \U26/Z_4 , \U26/Z_5 ,
         \U26/Z_6 , \U26/Z_7 , \U26/Z_8 , \U26/Z_9 , \U26/Z_10 , \U26/Z_11 ,
         \U26/Z_12 , \U26/Z_13 , \U26/Z_14 , \U26/Z_15 , \U26/Z_16 ,
         \U26/Z_17 , \U26/Z_18 , \U26/Z_19 , \U26/Z_20 , \U26/Z_21 ,
         \U26/Z_22 , \U26/Z_23 , \U26/Z_24 , \U26/Z_25 , \U26/Z_26 ,
         \U26/Z_27 , \U26/Z_28 , \U26/Z_29 , \U26/Z_30 , \U26/Z_31 ,
         \U26/Z_32 , \U26/Z_33 , \U26/Z_34 , \U26/Z_35 , \U26/Z_36 ,
         \U26/Z_37 , \U26/Z_38 , \U26/Z_39 , \U26/Z_40 , \U26/Z_41 ,
         \U26/Z_42 , \U26/Z_43 , \U26/Z_44 , \U26/Z_45 , \U26/Z_46 ,
         \U26/Z_47 , \U26/Z_48 , \U26/Z_49 , \U26/Z_50 , \U26/Z_51 ,
         \U26/Z_52 , \U26/Z_53 , \U26/Z_54 , \U26/Z_55 , \U26/Z_56 ,
         \U26/Z_57 , \U26/Z_58 , \U26/Z_59 , \U26/Z_60 , \U26/Z_61 ,
         \U26/Z_62 , \U26/Z_63 , \U26/Z_64 , \U26/Z_65 , \U26/Z_66 ,
         \U26/Z_67 , \U26/Z_68 , \U26/Z_69 , \U26/Z_70 , \U26/Z_71 ,
         \U26/Z_72 , \U26/Z_73 , \U26/Z_74 , \U26/Z_75 , \U26/Z_76 ,
         \U26/Z_77 , \U26/Z_78 , \U26/Z_79 , \U26/Z_80 , \U26/Z_81 ,
         \U26/Z_82 , \U26/Z_83 , \U26/Z_84 , \U26/Z_85 , \U26/Z_86 ,
         \U26/Z_87 , \U26/Z_88 , \U26/Z_89 , \U26/Z_90 , \U26/Z_91 ,
         \U26/Z_92 , \U26/Z_93 , \U26/Z_94 , \U26/Z_95 , \U26/Z_96 ,
         \U26/Z_97 , \U26/Z_98 , \U26/Z_99 , \U26/Z_100 , \U26/Z_101 ,
         \U26/Z_102 , \U26/Z_103 , \U26/Z_104 , \U26/Z_105 , \U26/Z_106 ,
         \U26/Z_107 , \U26/Z_108 , \U26/Z_109 , \U26/Z_110 , \U26/Z_111 ,
         \U26/Z_112 , \U26/Z_113 , \U26/Z_114 , \U26/Z_115 , \U26/Z_116 ,
         \U26/Z_117 , \U26/Z_118 , \U26/Z_119 , \U26/Z_120 , \U26/Z_121 ,
         \U26/Z_122 , \U26/Z_123 , \U26/Z_124 , \U26/Z_125 , \U26/Z_126 ,
         \U26/Z_127 , \U26/DATA1_0 , \U26/DATA1_1 , \U26/DATA1_2 ,
         \U26/DATA1_3 , \U26/DATA1_4 , \U26/DATA1_5 , \U26/DATA1_6 ,
         \U26/DATA1_7 , \U26/DATA1_8 , \U26/DATA1_9 , \U26/DATA1_10 ,
         \U26/DATA1_11 , \U26/DATA1_12 , \U26/DATA1_13 , \U26/DATA1_14 ,
         \U26/DATA1_15 , \U26/DATA1_16 , \U26/DATA1_17 , \U26/DATA1_18 ,
         \U26/DATA1_19 , \U26/DATA1_20 , \U26/DATA1_21 , \U26/DATA1_22 ,
         \U26/DATA1_23 , \U26/DATA1_24 , \U26/DATA1_25 , \U26/DATA1_26 ,
         \U26/DATA1_27 , \U26/DATA1_28 , \U26/DATA1_29 , \U26/DATA1_30 ,
         \U26/DATA1_31 , \U26/DATA1_32 , \U26/DATA1_33 , \U26/DATA1_34 ,
         \U26/DATA1_35 , \U26/DATA1_36 , \U26/DATA1_37 , \U26/DATA1_38 ,
         \U26/DATA1_39 , \U26/DATA1_40 , \U26/DATA1_41 , \U26/DATA1_42 ,
         \U26/DATA1_43 , \U26/DATA1_44 , \U26/DATA1_45 , \U26/DATA1_46 ,
         \U26/DATA1_47 , \U26/DATA1_48 , \U26/DATA1_49 , \U26/DATA1_50 ,
         \U26/DATA1_51 , \U26/DATA1_52 , \U26/DATA1_53 , \U26/DATA1_54 ,
         \U26/DATA1_55 , \U26/DATA1_56 , \U26/DATA1_57 , \U26/DATA1_58 ,
         \U26/DATA1_59 , \U26/DATA1_60 , \U26/DATA1_61 , \U26/DATA1_62 ,
         \U26/DATA1_63 , \U26/DATA1_64 , \U26/DATA1_65 , \U26/DATA1_66 ,
         \U26/DATA1_67 , \U26/DATA1_68 , \U26/DATA1_69 , \U26/DATA1_70 ,
         \U26/DATA1_71 , \U26/DATA1_72 , \U26/DATA1_73 , \U26/DATA1_74 ,
         \U26/DATA1_75 , \U26/DATA1_76 , \U26/DATA1_77 , \U26/DATA1_78 ,
         \U26/DATA1_79 , \U26/DATA1_80 , \U26/DATA1_81 , \U26/DATA1_82 ,
         \U26/DATA1_83 , \U26/DATA1_84 , \U26/DATA1_85 , \U26/DATA1_86 ,
         \U26/DATA1_87 , \U26/DATA1_88 , \U26/DATA1_89 , \U26/DATA1_90 ,
         \U26/DATA1_91 , \U26/DATA1_92 , \U26/DATA1_93 , \U26/DATA1_94 ,
         \U26/DATA1_95 , \U26/DATA1_96 , \U26/DATA1_97 , \U26/DATA1_98 ,
         \U26/DATA1_99 , \U26/DATA1_100 , \U26/DATA1_101 , \U26/DATA1_102 ,
         \U26/DATA1_103 , \U26/DATA1_104 , \U26/DATA1_105 , \U26/DATA1_106 ,
         \U26/DATA1_107 , \U26/DATA1_108 , \U26/DATA1_109 , \U26/DATA1_110 ,
         \U26/DATA1_111 , \U26/DATA1_112 , \U26/DATA1_113 , \U26/DATA1_114 ,
         \U26/DATA1_115 , \U26/DATA1_116 , \U26/DATA1_117 , \U26/DATA1_118 ,
         \U26/DATA1_119 , \U26/DATA1_120 , \U26/DATA1_121 , \U26/DATA1_122 ,
         \U26/DATA1_123 , \U26/DATA1_124 , \U26/DATA1_125 , \U26/DATA1_126 ,
         \U26/DATA1_127 , \U25/DATA2_0 , \U25/DATA2_1 , \U25/DATA2_2 ,
         \U25/DATA2_3 , \U25/DATA2_4 , \U25/DATA2_5 , \U25/DATA2_6 ,
         \U25/DATA2_7 , \U25/DATA2_8 , \U25/DATA2_9 , \U25/DATA2_10 ,
         \U25/DATA2_11 , \U25/DATA2_12 , \U25/DATA2_13 , \U25/DATA2_14 ,
         \U25/DATA2_15 , \U25/DATA2_16 , \U25/DATA2_17 , \U25/DATA2_18 ,
         \U25/DATA2_19 , \U25/DATA2_20 , \U25/DATA2_21 , \U25/DATA2_22 ,
         \U25/DATA2_23 , \U25/DATA2_24 , \U25/DATA2_25 , \U25/DATA2_26 ,
         \U25/DATA2_27 , \U25/DATA2_28 , \U25/DATA2_29 , \U25/DATA2_30 ,
         \U25/DATA2_31 , \U25/DATA2_32 , \U25/DATA2_33 , \U25/DATA2_34 ,
         \U25/DATA2_35 , \U24/Z_0 , \U24/DATA1_0 , \U23/Z_0 , \U23/DATA1_0 ,
         \U21/Z_0 , \U21/DATA1_0 , \U20/Z_0 , \U20/DATA1_0 , \U18/Z_0 ,
         \U18/Z_1 , \U18/Z_2 , \U18/Z_3 , \U18/Z_4 , \U18/Z_5 , \U18/Z_6 ,
         \U18/Z_7 , \U18/Z_8 , \U18/Z_9 , \U18/Z_10 , \U18/Z_11 , \U18/Z_12 ,
         \U18/Z_13 , \U18/Z_14 , \U18/Z_15 , \U18/Z_16 , \U18/Z_17 ,
         \U18/Z_18 , \U18/Z_19 , \U18/Z_20 , \U18/Z_21 , \U18/Z_22 ,
         \U18/Z_23 , \U18/Z_24 , \U18/Z_25 , \U18/Z_26 , \U18/Z_27 ,
         \U18/Z_28 , \U18/Z_29 , \U18/Z_30 , \U18/Z_31 , \U18/Z_32 ,
         \U18/Z_33 , \U18/Z_34 , \U18/Z_35 , \U17/Z_0 , \U17/DATA1_0 ,
         \U16/Z_0 , \U16/DATA1_0 , \U15/Z_0 , \U15/Z_1 , \U15/Z_2 , \U15/Z_3 ,
         \U15/Z_4 , \U15/Z_5 , \U15/Z_6 , \U15/Z_7 , \U15/DATA1_0 ,
         \U15/DATA1_1 , \U15/DATA1_2 , \U15/DATA1_3 , \U15/DATA1_4 ,
         \U15/DATA1_5 , \U15/DATA1_6 , \U15/DATA1_7 , \U14/Z_1 , \U14/Z_2 ,
         \U14/Z_3 , \U14/Z_4 , \U14/Z_5 , \U14/Z_6 , \U14/Z_7 , \U14/Z_8 ,
         \U14/Z_9 , \U14/Z_10 , \U14/Z_11 , \U14/Z_12 , \U14/Z_13 , \U14/Z_14 ,
         \U14/Z_15 , \U14/Z_16 , \U14/Z_17 , \U14/Z_18 , \U14/Z_19 ,
         \U14/Z_20 , \U14/Z_22 , \U14/Z_24 , \U14/Z_26 , \U14/Z_28 ,
         \U14/Z_30 , \U14/Z_32 , \U14/Z_34 , \U14/Z_35 , \U14/DATA1_21 ,
         \U14/DATA1_23 , \U14/DATA1_25 , \U14/DATA1_27 , \U14/DATA1_29 ,
         \U14/DATA1_31 , \U13/DATA1_3 , \U13/DATA1_4 , \U13/DATA1_5 ,
         \U13/DATA1_6 , \U12/Z_0 , \U5/DATA1_0 , \U5/DATA1_1 , \U5/DATA1_2 ,
         \U5/DATA1_3 , \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 , \U5/DATA1_7 ,
         \U5/DATA1_8 , \U5/DATA1_9 , \U5/DATA1_10 , \U5/DATA1_11 ,
         \U5/DATA1_12 , \U5/DATA1_13 , \U5/DATA1_14 , \U4/Z_3 , \U4/Z_4 ,
         \U4/Z_5 , \U4/Z_6 , n15, n18, n21, n24, n27, n30, n42, n43, n44, n45,
         n46, n47, n48, n49, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n157, n159, n165, n167, n171, n172,
         n209, n211, n212, n252, n253, n254, n255, n256, n257, n264, n265,
         n266, n269, n270, n271, n272, n273, n274, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n322, n323, n333, n337, n339, n340, n344, n345, n346, n350,
         n351, n352, n359, n362, n365, n368, n369, n371, n372, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n453, n454, n455, n456, n457, n458, n459,
         n510, n511, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1399,
         n1400, n1401, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977;
  assign \U36/DATA2_0  = m1ReadBus[0];
  assign \U36/DATA2_1  = m1ReadBus[1];
  assign \U36/DATA2_2  = m1ReadBus[2];
  assign \U36/DATA2_3  = m1ReadBus[3];
  assign \U36/DATA2_4  = m1ReadBus[4];
  assign \U36/DATA2_5  = m1ReadBus[5];
  assign \U36/DATA2_6  = m1ReadBus[6];
  assign \U36/DATA2_7  = m1ReadBus[7];
  assign \U36/DATA2_8  = m1ReadBus[8];
  assign \U36/DATA2_9  = m1ReadBus[9];
  assign \U36/DATA2_10  = m1ReadBus[10];
  assign \U36/DATA2_11  = m1ReadBus[11];
  assign \U36/DATA2_12  = m1ReadBus[12];
  assign \U36/DATA2_13  = m1ReadBus[13];
  assign \U36/DATA2_14  = m1ReadBus[14];
  assign \U36/DATA2_15  = m1ReadBus[15];
  assign \U36/DATA2_16  = m1ReadBus[16];
  assign \U36/DATA2_17  = m1ReadBus[17];
  assign \U36/DATA2_18  = m1ReadBus[18];
  assign \U36/DATA2_19  = m1ReadBus[19];
  assign \U36/DATA2_20  = m1ReadBus[20];
  assign \U36/DATA2_21  = m1ReadBus[21];
  assign \U36/DATA2_22  = m1ReadBus[22];
  assign \U36/DATA2_23  = m1ReadBus[23];
  assign \U36/DATA2_24  = m1ReadBus[24];
  assign \U36/DATA2_25  = m1ReadBus[25];
  assign \U36/DATA2_26  = m1ReadBus[26];
  assign \U36/DATA2_27  = m1ReadBus[27];
  assign \U36/DATA2_28  = m1ReadBus[28];
  assign \U36/DATA2_29  = m1ReadBus[29];
  assign \U36/DATA2_30  = m1ReadBus[30];
  assign \U36/DATA2_31  = m1ReadBus[31];
  assign \U36/DATA2_32  = m1ReadBus[32];
  assign \U36/DATA2_33  = m1ReadBus[33];
  assign \U36/DATA2_34  = m1ReadBus[34];
  assign \U36/DATA2_35  = m1ReadBus[35];
  assign \U36/DATA2_36  = m1ReadBus[36];
  assign \U36/DATA2_37  = m1ReadBus[37];
  assign \U36/DATA2_38  = m1ReadBus[38];
  assign \U36/DATA2_39  = m1ReadBus[39];
  assign \U36/DATA2_40  = m1ReadBus[40];
  assign \U36/DATA2_41  = m1ReadBus[41];
  assign \U36/DATA2_42  = m1ReadBus[42];
  assign \U36/DATA2_43  = m1ReadBus[43];
  assign \U36/DATA2_44  = m1ReadBus[44];
  assign \U36/DATA2_45  = m1ReadBus[45];
  assign \U36/DATA2_46  = m1ReadBus[46];
  assign \U36/DATA2_47  = m1ReadBus[47];
  assign \U36/DATA2_48  = m1ReadBus[48];
  assign \U36/DATA2_49  = m1ReadBus[49];
  assign \U36/DATA2_50  = m1ReadBus[50];
  assign \U36/DATA2_51  = m1ReadBus[51];
  assign \U36/DATA2_52  = m1ReadBus[52];
  assign \U36/DATA2_53  = m1ReadBus[53];
  assign \U36/DATA2_54  = m1ReadBus[54];
  assign \U36/DATA2_55  = m1ReadBus[55];
  assign \U36/DATA2_56  = m1ReadBus[56];
  assign \U36/DATA2_57  = m1ReadBus[57];
  assign \U36/DATA2_58  = m1ReadBus[58];
  assign \U36/DATA2_59  = m1ReadBus[59];
  assign \U36/DATA2_60  = m1ReadBus[60];
  assign \U36/DATA2_61  = m1ReadBus[61];
  assign \U36/DATA2_62  = m1ReadBus[62];
  assign \U36/DATA2_63  = m1ReadBus[63];
  assign \U36/DATA2_64  = m1ReadBus[64];
  assign \U36/DATA2_65  = m1ReadBus[65];
  assign \U36/DATA2_66  = m1ReadBus[66];
  assign \U36/DATA2_67  = m1ReadBus[67];
  assign \U36/DATA2_68  = m1ReadBus[68];
  assign \U36/DATA2_69  = m1ReadBus[69];
  assign \U36/DATA2_70  = m1ReadBus[70];
  assign \U36/DATA1_7  = m1ReadBus[71];
  assign \U36/DATA1_8  = m1ReadBus[72];
  assign \U36/DATA1_9  = m1ReadBus[73];
  assign \U36/DATA1_10  = m1ReadBus[74];
  assign \U36/DATA1_11  = m1ReadBus[75];
  assign \U36/DATA1_12  = m1ReadBus[76];
  assign \U36/DATA1_13  = m1ReadBus[77];
  assign \U36/DATA1_14  = m1ReadBus[78];
  assign \U36/DATA1_15  = m1ReadBus[79];
  assign \U36/DATA1_16  = m1ReadBus[80];
  assign \U36/DATA1_17  = m1ReadBus[81];
  assign \U36/DATA1_18  = m1ReadBus[82];
  assign \U36/DATA1_19  = m1ReadBus[83];
  assign \U36/DATA1_20  = m1ReadBus[84];
  assign \U36/DATA1_21  = m1ReadBus[85];
  assign \U36/DATA1_22  = m1ReadBus[86];
  assign \U36/DATA1_23  = m1ReadBus[87];
  assign \U36/DATA1_24  = m1ReadBus[88];
  assign \U36/DATA1_25  = m1ReadBus[89];
  assign \U36/DATA1_26  = m1ReadBus[90];
  assign \U36/DATA1_27  = m1ReadBus[91];
  assign \U36/DATA1_28  = m1ReadBus[92];
  assign \U36/DATA1_29  = m1ReadBus[93];
  assign \U36/DATA1_30  = m1ReadBus[94];
  assign \U36/DATA1_31  = m1ReadBus[95];
  assign \U36/DATA1_32  = m1ReadBus[96];
  assign \U36/DATA1_33  = m1ReadBus[97];
  assign \U36/DATA1_34  = m1ReadBus[98];
  assign \U36/DATA1_35  = m1ReadBus[99];
  assign \U36/DATA1_36  = m1ReadBus[100];
  assign \U36/DATA1_37  = m1ReadBus[101];
  assign \U36/DATA1_38  = m1ReadBus[102];
  assign \U36/DATA1_39  = m1ReadBus[103];
  assign \U36/DATA1_40  = m1ReadBus[104];
  assign \U36/DATA1_41  = m1ReadBus[105];
  assign \U36/DATA1_42  = m1ReadBus[106];
  assign \U36/DATA1_43  = m1ReadBus[107];
  assign \U36/DATA1_44  = m1ReadBus[108];
  assign \U36/DATA1_45  = m1ReadBus[109];
  assign \U36/DATA1_46  = m1ReadBus[110];
  assign \U36/DATA1_47  = m1ReadBus[111];
  assign \U36/DATA1_48  = m1ReadBus[112];
  assign \U36/DATA1_49  = m1ReadBus[113];
  assign \U36/DATA1_50  = m1ReadBus[114];
  assign \U36/DATA1_51  = m1ReadBus[115];
  assign \U36/DATA1_52  = m1ReadBus[116];
  assign \U36/DATA1_53  = m1ReadBus[117];
  assign \U36/DATA1_54  = m1ReadBus[118];
  assign \U36/DATA1_55  = m1ReadBus[119];
  assign \U36/DATA1_56  = m1ReadBus[120];
  assign \U36/DATA1_57  = m1ReadBus[121];
  assign \U36/DATA1_58  = m1ReadBus[122];
  assign \U36/DATA1_59  = m1ReadBus[123];
  assign \U36/DATA1_60  = m1ReadBus[124];
  assign \U36/DATA1_61  = m1ReadBus[125];
  assign \U36/DATA1_62  = m1ReadBus[126];
  assign \U36/DATA1_63  = m1ReadBus[127];
  assign m2ReadAddr[0] = \U29/Z_0 ;
  assign m2ReadAddr[1] = \U29/Z_1 ;
  assign m2ReadAddr[2] = \U29/Z_2 ;
  assign m2ReadAddr[3] = \U29/Z_3 ;
  assign m2ReadAddr[4] = \U29/Z_4 ;
  assign m2ReadAddr[5] = \U29/Z_5 ;
  assign m2ReadAddr[6] = \U29/Z_6 ;
  assign m2ReadAddr[7] = \U29/Z_7 ;
  assign m2WE = \U28/Z_0 ;
  assign m2WriteAddr[0] = \U27/Z_0 ;
  assign m2WriteAddr[1] = \U27/Z_1 ;
  assign m2WriteAddr[2] = \U27/Z_2 ;
  assign m2WriteAddr[3] = \U27/Z_3 ;
  assign m2WriteAddr[4] = \U27/Z_4 ;
  assign m2WriteAddr[5] = \U27/Z_5 ;
  assign m2WriteAddr[6] = \U27/Z_6 ;
  assign m2WriteAddr[7] = \U27/Z_7 ;
  assign m2WriteBus[0] = \U26/Z_0 ;
  assign m2WriteBus[1] = \U26/Z_1 ;
  assign m2WriteBus[2] = \U26/Z_2 ;
  assign m2WriteBus[3] = \U26/Z_3 ;
  assign m2WriteBus[4] = \U26/Z_4 ;
  assign m2WriteBus[5] = \U26/Z_5 ;
  assign m2WriteBus[6] = \U26/Z_6 ;
  assign m2WriteBus[7] = \U26/Z_7 ;
  assign m2WriteBus[8] = \U26/Z_8 ;
  assign m2WriteBus[9] = \U26/Z_9 ;
  assign m2WriteBus[10] = \U26/Z_10 ;
  assign m2WriteBus[11] = \U26/Z_11 ;
  assign m2WriteBus[12] = \U26/Z_12 ;
  assign m2WriteBus[13] = \U26/Z_13 ;
  assign m2WriteBus[14] = \U26/Z_14 ;
  assign m2WriteBus[15] = \U26/Z_15 ;
  assign m2WriteBus[16] = \U26/Z_16 ;
  assign m2WriteBus[17] = \U26/Z_17 ;
  assign m2WriteBus[18] = \U26/Z_18 ;
  assign m2WriteBus[19] = \U26/Z_19 ;
  assign m2WriteBus[20] = \U26/Z_20 ;
  assign m2WriteBus[21] = \U26/Z_21 ;
  assign m2WriteBus[22] = \U26/Z_22 ;
  assign m2WriteBus[23] = \U26/Z_23 ;
  assign m2WriteBus[24] = \U26/Z_24 ;
  assign m2WriteBus[25] = \U26/Z_25 ;
  assign m2WriteBus[26] = \U26/Z_26 ;
  assign m2WriteBus[27] = \U26/Z_27 ;
  assign m2WriteBus[28] = \U26/Z_28 ;
  assign m2WriteBus[29] = \U26/Z_29 ;
  assign m2WriteBus[30] = \U26/Z_30 ;
  assign m2WriteBus[31] = \U26/Z_31 ;
  assign m2WriteBus[32] = \U26/Z_32 ;
  assign m2WriteBus[33] = \U26/Z_33 ;
  assign m2WriteBus[34] = \U26/Z_34 ;
  assign m2WriteBus[35] = \U26/Z_35 ;
  assign m2WriteBus[36] = \U26/Z_36 ;
  assign m2WriteBus[37] = \U26/Z_37 ;
  assign m2WriteBus[38] = \U26/Z_38 ;
  assign m2WriteBus[39] = \U26/Z_39 ;
  assign m2WriteBus[40] = \U26/Z_40 ;
  assign m2WriteBus[41] = \U26/Z_41 ;
  assign m2WriteBus[42] = \U26/Z_42 ;
  assign m2WriteBus[43] = \U26/Z_43 ;
  assign m2WriteBus[44] = \U26/Z_44 ;
  assign m2WriteBus[45] = \U26/Z_45 ;
  assign m2WriteBus[46] = \U26/Z_46 ;
  assign m2WriteBus[47] = \U26/Z_47 ;
  assign m2WriteBus[48] = \U26/Z_48 ;
  assign m2WriteBus[49] = \U26/Z_49 ;
  assign m2WriteBus[50] = \U26/Z_50 ;
  assign m2WriteBus[51] = \U26/Z_51 ;
  assign m2WriteBus[52] = \U26/Z_52 ;
  assign m2WriteBus[53] = \U26/Z_53 ;
  assign m2WriteBus[54] = \U26/Z_54 ;
  assign m2WriteBus[55] = \U26/Z_55 ;
  assign m2WriteBus[56] = \U26/Z_56 ;
  assign m2WriteBus[57] = \U26/Z_57 ;
  assign m2WriteBus[58] = \U26/Z_58 ;
  assign m2WriteBus[59] = \U26/Z_59 ;
  assign m2WriteBus[60] = \U26/Z_60 ;
  assign m2WriteBus[61] = \U26/Z_61 ;
  assign m2WriteBus[62] = \U26/Z_62 ;
  assign m2WriteBus[63] = \U26/Z_63 ;
  assign m2WriteBus[64] = \U26/Z_64 ;
  assign m2WriteBus[65] = \U26/Z_65 ;
  assign m2WriteBus[66] = \U26/Z_66 ;
  assign m2WriteBus[67] = \U26/Z_67 ;
  assign m2WriteBus[68] = \U26/Z_68 ;
  assign m2WriteBus[69] = \U26/Z_69 ;
  assign m2WriteBus[70] = \U26/Z_70 ;
  assign m2WriteBus[71] = \U26/Z_71 ;
  assign m2WriteBus[72] = \U26/Z_72 ;
  assign m2WriteBus[73] = \U26/Z_73 ;
  assign m2WriteBus[74] = \U26/Z_74 ;
  assign m2WriteBus[75] = \U26/Z_75 ;
  assign m2WriteBus[76] = \U26/Z_76 ;
  assign m2WriteBus[77] = \U26/Z_77 ;
  assign m2WriteBus[78] = \U26/Z_78 ;
  assign m2WriteBus[79] = \U26/Z_79 ;
  assign m2WriteBus[80] = \U26/Z_80 ;
  assign m2WriteBus[81] = \U26/Z_81 ;
  assign m2WriteBus[82] = \U26/Z_82 ;
  assign m2WriteBus[83] = \U26/Z_83 ;
  assign m2WriteBus[84] = \U26/Z_84 ;
  assign m2WriteBus[85] = \U26/Z_85 ;
  assign m2WriteBus[86] = \U26/Z_86 ;
  assign m2WriteBus[87] = \U26/Z_87 ;
  assign m2WriteBus[88] = \U26/Z_88 ;
  assign m2WriteBus[89] = \U26/Z_89 ;
  assign m2WriteBus[90] = \U26/Z_90 ;
  assign m2WriteBus[91] = \U26/Z_91 ;
  assign m2WriteBus[92] = \U26/Z_92 ;
  assign m2WriteBus[93] = \U26/Z_93 ;
  assign m2WriteBus[94] = \U26/Z_94 ;
  assign m2WriteBus[95] = \U26/Z_95 ;
  assign m2WriteBus[96] = \U26/Z_96 ;
  assign m2WriteBus[97] = \U26/Z_97 ;
  assign m2WriteBus[98] = \U26/Z_98 ;
  assign m2WriteBus[99] = \U26/Z_99 ;
  assign m2WriteBus[100] = \U26/Z_100 ;
  assign m2WriteBus[101] = \U26/Z_101 ;
  assign m2WriteBus[102] = \U26/Z_102 ;
  assign m2WriteBus[103] = \U26/Z_103 ;
  assign m2WriteBus[104] = \U26/Z_104 ;
  assign m2WriteBus[105] = \U26/Z_105 ;
  assign m2WriteBus[106] = \U26/Z_106 ;
  assign m2WriteBus[107] = \U26/Z_107 ;
  assign m2WriteBus[108] = \U26/Z_108 ;
  assign m2WriteBus[109] = \U26/Z_109 ;
  assign m2WriteBus[110] = \U26/Z_110 ;
  assign m2WriteBus[111] = \U26/Z_111 ;
  assign m2WriteBus[112] = \U26/Z_112 ;
  assign m2WriteBus[113] = \U26/Z_113 ;
  assign m2WriteBus[114] = \U26/Z_114 ;
  assign m2WriteBus[115] = \U26/Z_115 ;
  assign m2WriteBus[116] = \U26/Z_116 ;
  assign m2WriteBus[117] = \U26/Z_117 ;
  assign m2WriteBus[118] = \U26/Z_118 ;
  assign m2WriteBus[119] = \U26/Z_119 ;
  assign m2WriteBus[120] = \U26/Z_120 ;
  assign m2WriteBus[121] = \U26/Z_121 ;
  assign m2WriteBus[122] = \U26/Z_122 ;
  assign m2WriteBus[123] = \U26/Z_123 ;
  assign m2WriteBus[124] = \U26/Z_124 ;
  assign m2WriteBus[125] = \U26/Z_125 ;
  assign m2WriteBus[126] = \U26/Z_126 ;
  assign m2WriteBus[127] = \U26/Z_127 ;
  assign \U25/DATA2_0  = m2ReadBus[0];
  assign \U25/DATA2_1  = m2ReadBus[1];
  assign \U25/DATA2_2  = m2ReadBus[2];
  assign \U25/DATA2_3  = m2ReadBus[3];
  assign \U25/DATA2_4  = m2ReadBus[4];
  assign \U25/DATA2_5  = m2ReadBus[5];
  assign \U25/DATA2_6  = m2ReadBus[6];
  assign \U25/DATA2_7  = m2ReadBus[7];
  assign \U25/DATA2_8  = m2ReadBus[8];
  assign \U25/DATA2_9  = m2ReadBus[9];
  assign \U25/DATA2_10  = m2ReadBus[10];
  assign \U25/DATA2_11  = m2ReadBus[11];
  assign \U25/DATA2_12  = m2ReadBus[12];
  assign \U25/DATA2_13  = m2ReadBus[13];
  assign \U25/DATA2_14  = m2ReadBus[14];
  assign \U25/DATA2_15  = m2ReadBus[15];
  assign \U25/DATA2_16  = m2ReadBus[16];
  assign \U25/DATA2_17  = m2ReadBus[17];
  assign \U25/DATA2_18  = m2ReadBus[18];
  assign \U25/DATA2_19  = m2ReadBus[19];
  assign \U25/DATA2_20  = m2ReadBus[20];
  assign \U25/DATA2_21  = m2ReadBus[21];
  assign \U25/DATA2_22  = m2ReadBus[22];
  assign \U25/DATA2_23  = m2ReadBus[23];
  assign \U25/DATA2_24  = m2ReadBus[24];
  assign \U25/DATA2_25  = m2ReadBus[25];
  assign \U25/DATA2_26  = m2ReadBus[26];
  assign \U25/DATA2_27  = m2ReadBus[27];
  assign \U25/DATA2_28  = m2ReadBus[28];
  assign \U25/DATA2_29  = m2ReadBus[29];
  assign \U25/DATA2_30  = m2ReadBus[30];
  assign \U25/DATA2_31  = m2ReadBus[31];
  assign \U25/DATA2_32  = m2ReadBus[32];
  assign \U25/DATA2_33  = m2ReadBus[33];
  assign \U25/DATA2_34  = m2ReadBus[34];
  assign \U25/DATA2_35  = m2ReadBus[35];
  assign m3WE = \U20/DATA1_0 ;
  assign m1ReadAddr[0] = \U5/DATA1_0 ;
  assign m1ReadAddr[1] = \U5/DATA1_1 ;
  assign m1ReadAddr[2] = \U5/DATA1_2 ;
  assign m1ReadAddr[3] = \U5/DATA1_3 ;
  assign m1ReadAddr[4] = \U5/DATA1_4 ;
  assign m1ReadAddr[5] = \U5/DATA1_5 ;
  assign m1ReadAddr[6] = \U5/DATA1_6 ;
  assign m1ReadAddr[7] = \U5/DATA1_7 ;
  assign m1ReadAddr[8] = \U5/DATA1_8 ;
  assign m1ReadAddr[9] = \U5/DATA1_9 ;
  assign m1ReadAddr[10] = \U5/DATA1_10 ;
  assign m1ReadAddr[11] = \U5/DATA1_11 ;
  assign m1ReadAddr[12] = \U5/DATA1_12 ;
  assign m1ReadAddr[13] = \U5/DATA1_13 ;
  assign m1ReadAddr[14] = \U5/DATA1_14 ;

  SDFFR_X2 write_enable_reg ( .D(1'b1), .SI(n211), .SE(n1368), .CK(clock), 
        .RN(n1636), .Q(\U23/DATA1_0 ) );
  SDFFR_X2 \readInitial_FS_reg[7]  ( .D(1'b0), .SI(n30), .SE(n1634), .CK(clock), .RN(n1636), .Q(\U15/DATA1_7 ), .QN(n1373) );
  SDFFR_X2 \readInitial_FS_reg[6]  ( .D(1'b0), .SI(n27), .SE(n1634), .CK(clock), .RN(n1636), .Q(\U15/DATA1_6 ), .QN(n1372) );
  SDFFR_X2 \readInitial_FS_reg[5]  ( .D(1'b0), .SI(n24), .SE(n1634), .CK(clock), .RN(n1636), .Q(\U15/DATA1_5 ) );
  SDFFR_X2 \readInitial_FS_reg[4]  ( .D(1'b0), .SI(n21), .SE(n1634), .CK(clock), .RN(n1636), .Q(\U15/DATA1_4 ) );
  SDFFR_X2 \readInitial_FS_reg[3]  ( .D(1'b0), .SI(n18), .SE(n1634), .CK(clock), .RN(n1636), .Q(\U15/DATA1_3 ) );
  SDFFR_X2 \readInitial_FS_reg[2]  ( .D(1'b0), .SI(n15), .SE(n1634), .CK(clock), .RN(n1636), .Q(\U15/DATA1_2 ) );
  SDFFR_X2 \readInitial_FS_reg[1]  ( .D(1'b0), .SI(\U29/DATA2_1 ), .SE(n1634), 
        .CK(clock), .RN(n1636), .Q(\U15/DATA1_1 ), .QN(n1374) );
  DFFS_X2 \scratchVal_FS_reg[21]  ( .D(\U18/Z_21 ), .CK(clock), .SN(n1636), 
        .Q(\U3/U1/DATA1_21 ) );
  DFFS_X2 \scratchVal_FS_reg[23]  ( .D(\U18/Z_23 ), .CK(clock), .SN(n1636), 
        .Q(\U3/U1/DATA1_23 ) );
  DFFS_X2 \scratchVal_FS_reg[25]  ( .D(\U18/Z_25 ), .CK(clock), .SN(n1636), 
        .Q(\U3/U1/DATA1_25 ) );
  DFFS_X2 \scratchVal_FS_reg[27]  ( .D(\U18/Z_27 ), .CK(clock), .SN(n1636), 
        .Q(\U3/U1/DATA1_27 ) );
  DFFS_X2 \scratchVal_FS_reg[29]  ( .D(\U18/Z_29 ), .CK(clock), .SN(n1636), 
        .Q(\U3/U1/DATA1_29 ) );
  DFFS_X2 \scratchVal_FS_reg[31]  ( .D(\U18/Z_31 ), .CK(clock), .SN(n1636), 
        .Q(\U3/U1/DATA1_31 ) );
  DFFS_X2 \scratchVal_FS_reg[33]  ( .D(\U18/Z_33 ), .CK(clock), .SN(rst_n), 
        .Q(\U3/U1/DATA1_33 ) );
  DFFS_X2 \scratchVal_Accum_reg[35]  ( .D(\U14/Z_35 ), .CK(clock), .SN(n1625), 
        .Q(\U3/U1/DATA2_35 ), .QN(n67) );
  DFFS_X2 \scratchVal_FS_reg[35]  ( .D(\U18/Z_35 ), .CK(clock), .SN(n1636), 
        .Q(\U3/U1/DATA1_35 ) );
  NAND2_X2 U162 ( .A1(\U29/DATA1_7 ), .A2(n1365), .ZN(n252) );
  NAND2_X2 U164 ( .A1(\U29/DATA1_6 ), .A2(n1623), .ZN(n253) );
  NAND2_X2 U166 ( .A1(\U29/DATA1_5 ), .A2(n1365), .ZN(n254) );
  NAND2_X2 U168 ( .A1(\U29/DATA1_4 ), .A2(n1623), .ZN(n255) );
  NAND2_X2 U170 ( .A1(\U29/DATA1_3 ), .A2(n1365), .ZN(n256) );
  NAND2_X2 U172 ( .A1(\U29/DATA1_2 ), .A2(n1623), .ZN(n257) );
  NAND2_X2 U186 ( .A1(\U29/DATA1_1 ), .A2(n1365), .ZN(n264) );
  NAND2_X2 U188 ( .A1(\U29/DATA1_0 ), .A2(n1623), .ZN(n265) );
  NAND2_X2 U190 ( .A1(\U28/DATA1_0 ), .A2(n1365), .ZN(n266) );
  NAND2_X2 U196 ( .A1(\U27/DATA1_7 ), .A2(n1623), .ZN(n269) );
  NAND2_X2 U198 ( .A1(\U27/DATA1_6 ), .A2(n1365), .ZN(n270) );
  NAND2_X2 U200 ( .A1(\U27/DATA1_5 ), .A2(n1623), .ZN(n271) );
  NAND2_X2 U202 ( .A1(\U27/DATA1_4 ), .A2(n1365), .ZN(n272) );
  NAND2_X2 U204 ( .A1(\U27/DATA1_3 ), .A2(n1623), .ZN(n273) );
  NAND2_X2 U206 ( .A1(\U27/DATA1_2 ), .A2(n1365), .ZN(n274) );
  NAND2_X2 U220 ( .A1(\U27/DATA1_1 ), .A2(n1365), .ZN(n281) );
  NAND2_X2 U222 ( .A1(\U27/DATA1_0 ), .A2(n1623), .ZN(n282) );
  NAND2_X2 U224 ( .A1(\U26/DATA1_9 ), .A2(n1365), .ZN(n283) );
  NAND2_X2 U226 ( .A1(\U26/DATA1_8 ), .A2(n1623), .ZN(n284) );
  NAND2_X2 U228 ( .A1(\U26/DATA1_7 ), .A2(n1365), .ZN(n285) );
  NAND2_X2 U230 ( .A1(\U26/DATA1_6 ), .A2(n1623), .ZN(n286) );
  NAND2_X2 U232 ( .A1(\U26/DATA1_5 ), .A2(n1365), .ZN(n287) );
  NAND2_X2 U234 ( .A1(\U26/DATA1_4 ), .A2(n1623), .ZN(n288) );
  NAND2_X2 U236 ( .A1(\U26/DATA1_35 ), .A2(n1365), .ZN(n289) );
  NAND2_X2 U238 ( .A1(\U26/DATA1_34 ), .A2(n1623), .ZN(n290) );
  NAND2_X2 U240 ( .A1(\U26/DATA1_33 ), .A2(n1365), .ZN(n291) );
  NAND2_X2 U242 ( .A1(\U26/DATA1_32 ), .A2(n1623), .ZN(n292) );
  NAND2_X2 U244 ( .A1(\U26/DATA1_31 ), .A2(n1365), .ZN(n293) );
  NAND2_X2 U246 ( .A1(\U26/DATA1_30 ), .A2(n1623), .ZN(n294) );
  NAND2_X2 U248 ( .A1(\U26/DATA1_3 ), .A2(n1365), .ZN(n295) );
  NAND2_X2 U250 ( .A1(\U26/DATA1_29 ), .A2(n1623), .ZN(n296) );
  NAND2_X2 U252 ( .A1(\U26/DATA1_28 ), .A2(n1365), .ZN(n297) );
  NAND2_X2 U254 ( .A1(\U26/DATA1_27 ), .A2(n1623), .ZN(n298) );
  NAND2_X2 U256 ( .A1(\U26/DATA1_26 ), .A2(n1623), .ZN(n299) );
  NAND2_X2 U258 ( .A1(\U26/DATA1_25 ), .A2(n1623), .ZN(n300) );
  NAND2_X2 U260 ( .A1(\U26/DATA1_24 ), .A2(n1623), .ZN(n301) );
  NAND2_X2 U262 ( .A1(\U26/DATA1_23 ), .A2(n1623), .ZN(n302) );
  NAND2_X2 U264 ( .A1(\U26/DATA1_22 ), .A2(n1623), .ZN(n303) );
  NAND2_X2 U266 ( .A1(\U26/DATA1_21 ), .A2(n1623), .ZN(n304) );
  NAND2_X2 U268 ( .A1(\U26/DATA1_20 ), .A2(n1623), .ZN(n305) );
  NAND2_X2 U270 ( .A1(\U26/DATA1_2 ), .A2(n1623), .ZN(n306) );
  NAND2_X2 U272 ( .A1(\U26/DATA1_19 ), .A2(n1623), .ZN(n307) );
  NAND2_X2 U274 ( .A1(\U26/DATA1_18 ), .A2(n1623), .ZN(n308) );
  NAND2_X2 U276 ( .A1(\U26/DATA1_17 ), .A2(n1623), .ZN(n309) );
  NAND2_X2 U278 ( .A1(\U26/DATA1_16 ), .A2(n1623), .ZN(n310) );
  NAND2_X2 U280 ( .A1(\U26/DATA1_15 ), .A2(n1623), .ZN(n311) );
  NAND2_X2 U282 ( .A1(\U26/DATA1_14 ), .A2(n1623), .ZN(n312) );
  NAND2_X2 U284 ( .A1(\U26/DATA1_13 ), .A2(n1623), .ZN(n313) );
  NAND2_X2 U286 ( .A1(\U26/DATA1_12 ), .A2(n1623), .ZN(n314) );
  NAND2_X2 U288 ( .A1(\U26/DATA1_11 ), .A2(n1623), .ZN(n315) );
  NAND2_X2 U290 ( .A1(\U26/DATA1_10 ), .A2(n1623), .ZN(n316) );
  NAND2_X2 U292 ( .A1(\U26/DATA1_1 ), .A2(n1623), .ZN(n317) );
  NAND2_X2 U294 ( .A1(\U26/DATA1_0 ), .A2(n1365), .ZN(n318) );
  AOI221_X2 U323 ( .B1(n1362), .B2(\U36/DATA2_34 ), .C1(n1361), .C2(
        \U36/DATA2_66 ), .A(n1973), .ZN(n371) );
  NAND2_X2 U325 ( .A1(n374), .A2(n375), .ZN(n351) );
  OAI22_X2 U328 ( .A1(n376), .A2(n165), .B1(\U13/DATA1_4 ), .B2(n377), .ZN(
        n352) );
  AOI221_X2 U329 ( .B1(\U36/DATA2_42 ), .B2(n1362), .C1(\U36/DATA1_10 ), .C2(
        n1361), .A(n1972), .ZN(n377) );
  AOI221_X2 U331 ( .B1(\U36/DATA2_58 ), .B2(n1362), .C1(\U36/DATA1_26 ), .C2(
        n1361), .A(n1971), .ZN(n376) );
  OAI22_X2 U334 ( .A1(n380), .A2(n165), .B1(\U13/DATA1_4 ), .B2(n381), .ZN(
        n322) );
  AOI221_X2 U335 ( .B1(\U36/DATA2_46 ), .B2(n1362), .C1(\U36/DATA1_14 ), .C2(
        n1361), .A(n1970), .ZN(n381) );
  AOI221_X2 U337 ( .B1(\U36/DATA2_62 ), .B2(n1362), .C1(\U36/DATA1_30 ), .C2(
        n1361), .A(n1969), .ZN(n380) );
  NAND2_X2 U339 ( .A1(n384), .A2(n385), .ZN(n323) );
  AOI221_X2 U342 ( .B1(\U36/DATA1_38 ), .B2(n1359), .C1(\U36/DATA2_6 ), .C2(
        n1358), .A(n1977), .ZN(n386) );
  AOI221_X2 U346 ( .B1(n1362), .B2(\U36/DATA2_32 ), .C1(n1361), .C2(
        \U36/DATA2_64 ), .A(n1968), .ZN(n389) );
  OAI22_X2 U350 ( .A1(n394), .A2(n165), .B1(\U13/DATA1_4 ), .B2(n395), .ZN(
        n393) );
  AOI221_X2 U351 ( .B1(\U36/DATA2_40 ), .B2(n1362), .C1(\U36/DATA1_8 ), .C2(
        n1361), .A(n1967), .ZN(n395) );
  AOI221_X2 U353 ( .B1(\U36/DATA2_56 ), .B2(n1362), .C1(\U36/DATA1_24 ), .C2(
        n1361), .A(n1966), .ZN(n394) );
  OAI22_X2 U356 ( .A1(n398), .A2(n165), .B1(\U13/DATA1_4 ), .B2(n399), .ZN(
        n337) );
  AOI221_X2 U357 ( .B1(\U36/DATA2_44 ), .B2(n1362), .C1(\U36/DATA1_12 ), .C2(
        n1361), .A(n1965), .ZN(n399) );
  AOI221_X2 U359 ( .B1(\U36/DATA2_60 ), .B2(n1362), .C1(\U36/DATA1_28 ), .C2(
        n1361), .A(n1964), .ZN(n398) );
  NAND2_X2 U361 ( .A1(n402), .A2(n403), .ZN(n339) );
  AOI221_X2 U364 ( .B1(\U36/DATA1_36 ), .B2(n1359), .C1(\U36/DATA2_4 ), .C2(
        n1358), .A(n1976), .ZN(n404) );
  OAI22_X2 U369 ( .A1(n410), .A2(n165), .B1(\U13/DATA1_4 ), .B2(n411), .ZN(
        n409) );
  AOI221_X2 U370 ( .B1(\U36/DATA2_45 ), .B2(n1362), .C1(\U36/DATA1_13 ), .C2(
        n1361), .A(n1963), .ZN(n411) );
  AOI221_X2 U372 ( .B1(\U36/DATA2_61 ), .B2(n1362), .C1(\U36/DATA1_29 ), .C2(
        n1361), .A(n1962), .ZN(n410) );
  AOI221_X2 U376 ( .B1(\U36/DATA1_37 ), .B2(n1359), .C1(\U36/DATA2_5 ), .C2(
        n1358), .A(n1975), .ZN(n408) );
  OAI22_X2 U379 ( .A1(n419), .A2(n165), .B1(\U13/DATA1_4 ), .B2(n420), .ZN(
        n418) );
  AOI221_X2 U380 ( .B1(\U36/DATA2_41 ), .B2(n1362), .C1(\U36/DATA1_9 ), .C2(
        n1361), .A(n1961), .ZN(n420) );
  AOI221_X2 U382 ( .B1(\U36/DATA2_57 ), .B2(n1362), .C1(\U36/DATA1_25 ), .C2(
        n1361), .A(n1960), .ZN(n419) );
  AOI221_X2 U386 ( .B1(\U36/DATA1_33 ), .B2(n1359), .C1(\U36/DATA2_1 ), .C2(
        n1358), .A(n1974), .ZN(n417) );
  AOI221_X2 U390 ( .B1(n1362), .B2(\U36/DATA2_35 ), .C1(n1361), .C2(
        \U36/DATA2_67 ), .A(n1959), .ZN(n427) );
  NAND2_X2 U393 ( .A1(n429), .A2(n430), .ZN(n346) );
  NOR2_X2 U396 ( .A1(n165), .A2(\U13/DATA1_3 ), .ZN(n369) );
  OAI22_X2 U397 ( .A1(n431), .A2(n165), .B1(\U13/DATA1_4 ), .B2(n432), .ZN(
        n345) );
  AOI221_X2 U398 ( .B1(\U36/DATA2_43 ), .B2(n1362), .C1(\U36/DATA1_11 ), .C2(
        n1361), .A(n1958), .ZN(n432) );
  AOI221_X2 U400 ( .B1(\U36/DATA2_59 ), .B2(n1362), .C1(\U36/DATA1_27 ), .C2(
        n1361), .A(n1957), .ZN(n431) );
  NOR3_X2 U456 ( .A1(n457), .A2(n458), .A3(n459), .ZN(n456) );
  NAND2_X2 U457 ( .A1(\U25/DATA2_27 ), .A2(\U25/DATA2_25 ), .ZN(n459) );
  NAND3_X2 U458 ( .A1(\U25/DATA2_21 ), .A2(n1634), .A3(\U25/DATA2_23 ), .ZN(
        n458) );
  NAND4_X2 U459 ( .A1(\U25/DATA2_35 ), .A2(\U25/DATA2_33 ), .A3(\U25/DATA2_31 ), .A4(\U25/DATA2_29 ), .ZN(n457) );
  NOR4_X2 U460 ( .A1(\U25/DATA2_24 ), .A2(\U25/DATA2_22 ), .A3(\U25/DATA2_20 ), 
        .A4(n1462), .ZN(n455) );
  NOR3_X2 U461 ( .A1(\U25/DATA2_30 ), .A2(\U25/DATA2_34 ), .A3(\U25/DATA2_32 ), 
        .ZN(n454) );
  NOR2_X2 U462 ( .A1(\U25/DATA2_28 ), .A2(\U25/DATA2_26 ), .ZN(n453) );
  NAND2_X2 U513 ( .A1(n1368), .A2(n209), .ZN(\U12/Z_0 ) );
  NOR2_X2 U523 ( .A1(n165), .A2(n167), .ZN(n340) );
  AND2_X1 U699 ( .A1(\U24/DATA1_0 ), .A2(start), .ZN(\U24/Z_0 ) );
  AND2_X1 U700 ( .A1(\U23/DATA1_0 ), .A2(start), .ZN(\U23/Z_0 ) );
  AND2_X1 U701 ( .A1(n391), .A2(n392), .ZN(n365) );
  AND2_X1 U702 ( .A1(n414), .A2(n415), .ZN(n333) );
  AND2_X1 U703 ( .A1(n423), .A2(n424), .ZN(n359) );
  AND2_X1 U705 ( .A1(\U21/DATA1_0 ), .A2(start), .ZN(\U21/Z_0 ) );
  AND2_X1 U706 ( .A1(\U20/DATA1_0 ), .A2(start), .ZN(\U20/Z_0 ) );
  AND2_X1 U708 ( .A1(\U17/DATA1_0 ), .A2(start), .ZN(\U17/Z_0 ) );
  Cdf_top dut_CDF_top ( .clock(clock), .reset_n(n1624), .start(n1623), 
        .SP_ReadBus({m2ReadBus[127:36], \U25/DATA2_35 , \U25/DATA2_34 , 
        \U25/DATA2_33 , \U25/DATA2_32 , \U25/DATA2_31 , \U25/DATA2_30 , 
        \U25/DATA2_29 , \U25/DATA2_28 , \U25/DATA2_27 , \U25/DATA2_26 , 
        \U25/DATA2_25 , \U25/DATA2_24 , \U25/DATA2_23 , \U25/DATA2_22 , 
        \U25/DATA2_21 , \U25/DATA2_20 , \U25/DATA2_19 , \U25/DATA2_18 , 
        \U25/DATA2_17 , \U25/DATA2_16 , \U25/DATA2_15 , \U25/DATA2_14 , 
        \U25/DATA2_13 , \U25/DATA2_12 , \U25/DATA2_11 , \U25/DATA2_10 , 
        \U25/DATA2_9 , \U25/DATA2_8 , \U25/DATA2_7 , \U25/DATA2_6 , 
        \U25/DATA2_5 , \U25/DATA2_4 , \U25/DATA2_3 , \U25/DATA2_2 , 
        \U25/DATA2_1 , \U25/DATA2_0 }), .SP_ReadAddress({\U29/DATA1_15 , 
        \U29/DATA1_14 , \U29/DATA1_13 , \U29/DATA1_12 , \U29/DATA1_11 , 
        \U29/DATA1_10 , \U29/DATA1_9 , \U29/DATA1_8 , \U29/DATA1_7 , 
        \U29/DATA1_6 , \U29/DATA1_5 , \U29/DATA1_4 , \U29/DATA1_3 , 
        \U29/DATA1_2 , \U29/DATA1_1 , \U29/DATA1_0 }), .WriteEnable(
        \U28/DATA1_0 ), .Output_MEMBus({\U26/DATA1_127 , \U26/DATA1_126 , 
        \U26/DATA1_125 , \U26/DATA1_124 , \U26/DATA1_123 , \U26/DATA1_122 , 
        \U26/DATA1_121 , \U26/DATA1_120 , \U26/DATA1_119 , \U26/DATA1_118 , 
        \U26/DATA1_117 , \U26/DATA1_116 , \U26/DATA1_115 , \U26/DATA1_114 , 
        \U26/DATA1_113 , \U26/DATA1_112 , \U26/DATA1_111 , \U26/DATA1_110 , 
        \U26/DATA1_109 , \U26/DATA1_108 , \U26/DATA1_107 , \U26/DATA1_106 , 
        \U26/DATA1_105 , \U26/DATA1_104 , \U26/DATA1_103 , \U26/DATA1_102 , 
        \U26/DATA1_101 , \U26/DATA1_100 , \U26/DATA1_99 , \U26/DATA1_98 , 
        \U26/DATA1_97 , \U26/DATA1_96 , \U26/DATA1_95 , \U26/DATA1_94 , 
        \U26/DATA1_93 , \U26/DATA1_92 , \U26/DATA1_91 , \U26/DATA1_90 , 
        \U26/DATA1_89 , \U26/DATA1_88 , \U26/DATA1_87 , \U26/DATA1_86 , 
        \U26/DATA1_85 , \U26/DATA1_84 , \U26/DATA1_83 , \U26/DATA1_82 , 
        \U26/DATA1_81 , \U26/DATA1_80 , \U26/DATA1_79 , \U26/DATA1_78 , 
        \U26/DATA1_77 , \U26/DATA1_76 , \U26/DATA1_75 , \U26/DATA1_74 , 
        \U26/DATA1_73 , \U26/DATA1_72 , \U26/DATA1_71 , \U26/DATA1_70 , 
        \U26/DATA1_69 , \U26/DATA1_68 , \U26/DATA1_67 , \U26/DATA1_66 , 
        \U26/DATA1_65 , \U26/DATA1_64 , \U26/DATA1_63 , \U26/DATA1_62 , 
        \U26/DATA1_61 , \U26/DATA1_60 , \U26/DATA1_59 , \U26/DATA1_58 , 
        \U26/DATA1_57 , \U26/DATA1_56 , \U26/DATA1_55 , \U26/DATA1_54 , 
        \U26/DATA1_53 , \U26/DATA1_52 , \U26/DATA1_51 , \U26/DATA1_50 , 
        \U26/DATA1_49 , \U26/DATA1_48 , \U26/DATA1_47 , \U26/DATA1_46 , 
        \U26/DATA1_45 , \U26/DATA1_44 , \U26/DATA1_43 , \U26/DATA1_42 , 
        \U26/DATA1_41 , \U26/DATA1_40 , \U26/DATA1_39 , \U26/DATA1_38 , 
        \U26/DATA1_37 , \U26/DATA1_36 , \U26/DATA1_35 , \U26/DATA1_34 , 
        \U26/DATA1_33 , \U26/DATA1_32 , \U26/DATA1_31 , \U26/DATA1_30 , 
        \U26/DATA1_29 , \U26/DATA1_28 , \U26/DATA1_27 , \U26/DATA1_26 , 
        \U26/DATA1_25 , \U26/DATA1_24 , \U26/DATA1_23 , \U26/DATA1_22 , 
        \U26/DATA1_21 , \U26/DATA1_20 , \U26/DATA1_19 , \U26/DATA1_18 , 
        \U26/DATA1_17 , \U26/DATA1_16 , \U26/DATA1_15 , \U26/DATA1_14 , 
        \U26/DATA1_13 , \U26/DATA1_12 , \U26/DATA1_11 , \U26/DATA1_10 , 
        \U26/DATA1_9 , \U26/DATA1_8 , \U26/DATA1_7 , \U26/DATA1_6 , 
        \U26/DATA1_5 , \U26/DATA1_4 , \U26/DATA1_3 , \U26/DATA1_2 , 
        \U26/DATA1_1 , \U26/DATA1_0 }), .Output_MEMAddress({\U27/DATA1_15 , 
        \U27/DATA1_14 , \U27/DATA1_13 , \U27/DATA1_12 , \U27/DATA1_11 , 
        \U27/DATA1_10 , \U27/DATA1_9 , \U27/DATA1_8 , \U27/DATA1_7 , 
        \U27/DATA1_6 , \U27/DATA1_5 , \U27/DATA1_4 , \U27/DATA1_3 , 
        \U27/DATA1_2 , \U27/DATA1_1 , \U27/DATA1_0 }), .Cdf_Min(cdf_min), 
        .done(done), .input_base_offset(inputBaseOffset), .cdf_valid(cdf_valid) );
  DFFR_X2 \pipelineCounter_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .RN(n1624), .Q(
        \U13/DATA1_3 ), .QN(n167) );
  DFFR_X2 \pipelineCounter_reg[4]  ( .D(\U4/Z_4 ), .CK(clock), .RN(n1624), .Q(
        \U13/DATA1_4 ), .QN(n165) );
  DFFS_X2 \scratchVal_Accum_reg[25]  ( .D(n1471), .CK(clock), .SN(rst_n), .Q(
        n1811), .QN(n77) );
  DFFS_X2 \scratchVal_Accum_reg[33]  ( .D(n1470), .CK(clock), .SN(n1624), .Q(
        n1860), .QN(n69) );
  DFFS_X2 \scratchVal_Accum_reg[27]  ( .D(n1469), .CK(clock), .SN(n1625), .Q(
        n1825), .QN(n75) );
  DFFR_X2 \readInitial_Accum_reg[3]  ( .D(\U15/Z_3 ), .CK(clock), .RN(n1624), 
        .Q(\U27/DATA2_3 ), .QN(n46) );
  DFFR_X2 \readInitial_Accum_reg[1]  ( .D(\U15/Z_1 ), .CK(clock), .RN(n1624), 
        .Q(\U27/DATA2_1 ), .QN(n48) );
  DFFR_X2 \memoryCounter_reg[14]  ( .D(n510), .CK(clock), .RN(n1625), .Q(
        \U5/DATA1_14 ), .QN(n171) );
  SDFFS_X2 \scratchVal_Accum_reg[31]  ( .D(n1635), .SI(1'b1), .SE(
        \U14/DATA1_31 ), .CK(clock), .SN(n1626), .Q(n1364), .QN(n71) );
  DFFR_X2 \memoryCounter_reg[13]  ( .D(n1955), .CK(clock), .RN(n1626), .Q(
        \U5/DATA1_13 ), .QN(n1463) );
  DFFR_X2 \readInitial_Accum_reg[2]  ( .D(\U15/Z_2 ), .CK(clock), .RN(n1624), 
        .Q(\U27/DATA2_2 ), .QN(n47) );
  DFFR_X2 \memoryCounter_reg[0]  ( .D(n511), .CK(clock), .RN(n1636), .Q(
        \U5/DATA1_0 ), .QN(n172) );
  DFFR_X2 \readInitial_Accum_reg[4]  ( .D(\U15/Z_4 ), .CK(clock), .RN(n1624), 
        .Q(\U27/DATA2_4 ), .QN(n45) );
  DFFR_X2 \scratchVal_Accum_reg[0]  ( .D(n1403), .CK(clock), .RN(rst_n), .Q(
        n1673), .QN(n102) );
  SDFFR_X1 \readInitial_FS_reg[0]  ( .D(1'b0), .SI(\U29/DATA2_0 ), .SE(start), 
        .CK(clock), .RN(rst_n), .Q(\U15/DATA1_0 ), .QN(n1646) );
  DFFS_X2 \scratchVal_Accum_reg[23]  ( .D(n1401), .CK(clock), .SN(rst_n), .Q(
        n1804), .QN(n79) );
  DFFS_X2 \scratchVal_Accum_reg[29]  ( .D(n1400), .CK(clock), .SN(n1636), .Q(
        n1844), .QN(n73) );
  DFFS_X2 \scratchVal_Accum_reg[21]  ( .D(n1399), .CK(clock), .SN(n1636), .Q(
        n1796), .QN(n81) );
  SDFFR_X1 \readInitial_FI_reg[7]  ( .D(n1634), .SI(1'b0), .SE(n344), .CK(
        clock), .RN(n1636), .Q(n30), .QN(n59) );
  SDFFR_X1 \readInitial_FI_reg[5]  ( .D(1'b0), .SI(n1634), .SE(n1640), .CK(
        clock), .RN(n1636), .Q(n24), .QN(n61) );
  SDFFR_X1 \readInitial_FI_reg[1]  ( .D(1'b0), .SI(n1634), .SE(n1649), .CK(
        clock), .RN(n1636), .Q(\U29/DATA2_1 ), .QN(n65) );
  SDFFR_X1 \readInitial_FI_reg[0]  ( .D(1'b0), .SI(n1634), .SE(n1645), .CK(
        clock), .RN(n1636), .Q(\U29/DATA2_0 ), .QN(n66) );
  SDFFR_X1 \readInitial_FI_reg[3]  ( .D(n1634), .SI(1'b0), .SE(n426), .CK(
        clock), .RN(n1636), .Q(n18), .QN(n63) );
  SDFFR_X1 \readInitial_FI_reg[2]  ( .D(n1634), .SI(1'b0), .SE(n368), .CK(
        clock), .RN(n1636), .Q(n15), .QN(n64) );
  SDFFR_X1 \readInitial_FI_reg[6]  ( .D(n1634), .SI(1'b0), .SE(n350), .CK(
        clock), .RN(n1636), .Q(n27), .QN(n60) );
  SDFFR_X1 \readInitial_FI_reg[4]  ( .D(n1634), .SI(1'b0), .SE(n362), .CK(
        clock), .RN(n1636), .Q(n21), .QN(n62) );
  DFFR_X2 m2WE_Accum_reg ( .D(\U16/Z_0 ), .CK(clock), .RN(n1625), .Q(n1366), 
        .QN(n1665) );
  DFFR_X2 \readInitial_Accum_reg[7]  ( .D(\U15/Z_7 ), .CK(clock), .RN(n1624), 
        .Q(\U27/DATA2_7 ), .QN(n42) );
  DFFR_X2 \readInitial_Accum_reg[6]  ( .D(\U15/Z_6 ), .CK(clock), .RN(n1624), 
        .Q(\U27/DATA2_6 ), .QN(n43) );
  DFFR_X2 \readInitial_Accum_reg[5]  ( .D(\U15/Z_5 ), .CK(clock), .RN(n1624), 
        .Q(\U27/DATA2_5 ), .QN(n44) );
  DFFR_X2 \readInitial_Accum_reg[0]  ( .D(\U15/Z_0 ), .CK(clock), .RN(n1636), 
        .Q(\U27/DATA2_0 ), .QN(n49) );
  DFFR_X2 \pipelineCounter_reg[6]  ( .D(\U4/Z_6 ), .CK(clock), .RN(n1625), .Q(
        \U13/DATA1_6 ), .QN(n157) );
  DFFR_X2 \pipelineCounter_reg[5]  ( .D(\U4/Z_5 ), .CK(clock), .RN(n1626), .Q(
        \U13/DATA1_5 ), .QN(n159) );
  DFFR_X2 \scratchVal_Accum_reg[1]  ( .D(\U14/Z_1 ), .CK(clock), .RN(n1636), 
        .Q(n1677), .QN(n101) );
  DFFR_X2 \scratchVal_Accum_reg[2]  ( .D(\U14/Z_2 ), .CK(clock), .RN(n1636), 
        .Q(n1681), .QN(n100) );
  DFFR_X2 \scratchVal_Accum_reg[3]  ( .D(\U14/Z_3 ), .CK(clock), .RN(n1636), 
        .Q(n1686), .QN(n99) );
  DFFR_X2 \scratchVal_Accum_reg[9]  ( .D(\U14/Z_9 ), .CK(clock), .RN(n1636), 
        .Q(n1721), .QN(n93) );
  DFFR_X2 \scratchVal_Accum_reg[4]  ( .D(\U14/Z_4 ), .CK(clock), .RN(n1636), 
        .Q(n1690), .QN(n98) );
  DFFR_X2 \scratchVal_Accum_reg[10]  ( .D(\U14/Z_10 ), .CK(clock), .RN(n1636), 
        .Q(n1725), .QN(n92) );
  DFFR_X2 \scratchVal_Accum_reg[5]  ( .D(\U14/Z_5 ), .CK(clock), .RN(n1636), 
        .Q(n1695), .QN(n97) );
  DFFR_X2 \scratchVal_Accum_reg[15]  ( .D(\U14/Z_15 ), .CK(clock), .RN(n1636), 
        .Q(n1756), .QN(n87) );
  DFFR_X2 \scratchVal_Accum_reg[11]  ( .D(\U14/Z_11 ), .CK(clock), .RN(n1636), 
        .Q(n1729), .QN(n91) );
  DFFR_X2 \scratchVal_Accum_reg[30]  ( .D(\U14/Z_30 ), .CK(clock), .RN(n1636), 
        .Q(n1849), .QN(n72) );
  DFFR_X2 \scratchVal_Accum_reg[22]  ( .D(\U14/Z_22 ), .CK(clock), .RN(n1636), 
        .Q(n1802), .QN(n80) );
  DFFR_X2 \scratchVal_Accum_reg[16]  ( .D(\U14/Z_16 ), .CK(clock), .RN(n1636), 
        .Q(n1760), .QN(n86) );
  DFFR_X2 \scratchVal_Accum_reg[6]  ( .D(\U14/Z_6 ), .CK(clock), .RN(rst_n), 
        .Q(n1699), .QN(n96) );
  DFFR_X2 \scratchVal_Accum_reg[24]  ( .D(\U14/Z_24 ), .CK(clock), .RN(n1636), 
        .Q(n1808), .QN(n78) );
  DFFR_X2 \scratchVal_Accum_reg[12]  ( .D(\U14/Z_12 ), .CK(clock), .RN(n1636), 
        .Q(n1733), .QN(n90) );
  DFFR_X2 \scratchVal_Accum_reg[7]  ( .D(\U14/Z_7 ), .CK(clock), .RN(n1636), 
        .Q(n1703), .QN(n95) );
  DFFR_X2 \scratchVal_Accum_reg[32]  ( .D(\U14/Z_32 ), .CK(clock), .RN(rst_n), 
        .Q(n1857), .QN(n70) );
  DFFR_X2 \scratchVal_Accum_reg[8]  ( .D(\U14/Z_8 ), .CK(clock), .RN(n1636), 
        .Q(n1709), .QN(n94) );
  DFFR_X2 \scratchVal_Accum_reg[19]  ( .D(\U14/Z_19 ), .CK(clock), .RN(n1624), 
        .Q(n1775), .QN(n83) );
  DFFR_X2 \scratchVal_Accum_reg[13]  ( .D(\U14/Z_13 ), .CK(clock), .RN(n1636), 
        .Q(n1737), .QN(n89) );
  DFFR_X2 \scratchVal_Accum_reg[17]  ( .D(\U14/Z_17 ), .CK(clock), .RN(n1625), 
        .Q(n1765), .QN(n85) );
  DFFR_X2 \scratchVal_Accum_reg[20]  ( .D(\U14/Z_20 ), .CK(clock), .RN(n1626), 
        .Q(n1779), .QN(n82) );
  DFFR_X2 \scratchVal_Accum_reg[18]  ( .D(\U14/Z_18 ), .CK(clock), .RN(rst_n), 
        .Q(n1769), .QN(n84) );
  DFFR_X2 \scratchVal_Accum_reg[34]  ( .D(\U14/Z_34 ), .CK(clock), .RN(n1624), 
        .Q(n1867), .QN(n68) );
  DFFR_X2 \scratchVal_Accum_reg[14]  ( .D(\U14/Z_14 ), .CK(clock), .RN(n1636), 
        .Q(n1744), .QN(n88) );
  DFFR_X2 \scratchVal_Accum_reg[28]  ( .D(\U14/Z_28 ), .CK(clock), .RN(n1625), 
        .Q(n1832), .QN(n74) );
  DFFR_X2 \scratchVal_Accum_reg[26]  ( .D(\U14/Z_26 ), .CK(clock), .RN(n1626), 
        .Q(n1816), .QN(n76) );
  DFFR_X2 m2WE_FS_reg ( .D(\U20/Z_0 ), .CK(clock), .RN(n1626), .Q(
        \U16/DATA1_0 ) );
  DFFR_X2 m2WE_FI_reg ( .D(\U23/Z_0 ), .CK(clock), .RN(n1625), .Q(
        \U20/DATA1_0 ) );
  DFFR_X2 done_FS_reg ( .D(\U21/Z_0 ), .CK(clock), .RN(n1626), .Q(
        \U17/DATA1_0 ) );
  DFFR_X2 done_FI_reg ( .D(\U24/Z_0 ), .CK(clock), .RN(n1625), .Q(
        \U21/DATA1_0 ) );
  DFFR_X2 done_Accum_reg ( .D(\U17/Z_0 ), .CK(clock), .RN(n1625), .Q(n1365), 
        .QN(n1633) );
  DFFR_X2 \scratchVal_FS_reg[34]  ( .D(\U18/Z_34 ), .CK(clock), .RN(rst_n), 
        .Q(\U3/U1/DATA1_34 ) );
  DFFR_X2 \scratchVal_FS_reg[32]  ( .D(\U18/Z_32 ), .CK(clock), .RN(n1624), 
        .Q(\U3/U1/DATA1_32 ) );
  DFFR_X2 \scratchVal_FS_reg[30]  ( .D(\U18/Z_30 ), .CK(clock), .RN(n1626), 
        .Q(\U3/U1/DATA1_30 ) );
  DFFR_X2 \scratchVal_FS_reg[28]  ( .D(\U18/Z_28 ), .CK(clock), .RN(rst_n), 
        .Q(\U3/U1/DATA1_28 ) );
  DFFR_X2 \scratchVal_FS_reg[26]  ( .D(\U18/Z_26 ), .CK(clock), .RN(n1624), 
        .Q(\U3/U1/DATA1_26 ) );
  DFFR_X2 \scratchVal_FS_reg[24]  ( .D(\U18/Z_24 ), .CK(clock), .RN(rst_n), 
        .Q(\U3/U1/DATA1_24 ) );
  DFFR_X2 \scratchVal_FS_reg[22]  ( .D(\U18/Z_22 ), .CK(clock), .RN(n1624), 
        .Q(\U3/U1/DATA1_22 ) );
  DFFR_X2 \scratchVal_FS_reg[20]  ( .D(\U18/Z_20 ), .CK(clock), .RN(rst_n), 
        .Q(\U3/U1/DATA1_20 ) );
  DFFR_X2 done_enable_reg ( .D(n1956), .CK(clock), .RN(n1626), .Q(
        \U24/DATA1_0 ) );
  DFFR_X2 \scratchVal_FS_reg[19]  ( .D(\U18/Z_19 ), .CK(clock), .RN(rst_n), 
        .Q(\U3/U1/DATA1_19 ) );
  DFFR_X2 \scratchVal_FS_reg[18]  ( .D(\U18/Z_18 ), .CK(clock), .RN(rst_n), 
        .Q(\U3/U1/DATA1_18 ) );
  DFFR_X2 \scratchVal_FS_reg[17]  ( .D(\U18/Z_17 ), .CK(clock), .RN(rst_n), 
        .Q(\U3/U1/DATA1_17 ) );
  DFFR_X2 \scratchVal_FS_reg[16]  ( .D(\U18/Z_16 ), .CK(clock), .RN(n1636), 
        .Q(\U3/U1/DATA1_16 ) );
  DFFR_X2 \scratchVal_FS_reg[15]  ( .D(\U18/Z_15 ), .CK(clock), .RN(n1636), 
        .Q(\U3/U1/DATA1_15 ) );
  DFFR_X2 \scratchVal_FS_reg[14]  ( .D(\U18/Z_14 ), .CK(clock), .RN(n1636), 
        .Q(\U3/U1/DATA1_14 ) );
  DFFR_X2 \scratchVal_FS_reg[13]  ( .D(\U18/Z_13 ), .CK(clock), .RN(n1636), 
        .Q(\U3/U1/DATA1_13 ) );
  DFFR_X2 \scratchVal_FS_reg[12]  ( .D(\U18/Z_12 ), .CK(clock), .RN(n1636), 
        .Q(\U3/U1/DATA1_12 ) );
  DFFR_X2 \scratchVal_FS_reg[11]  ( .D(\U18/Z_11 ), .CK(clock), .RN(n1636), 
        .Q(\U3/U1/DATA1_11 ) );
  DFFR_X2 \scratchVal_FS_reg[10]  ( .D(\U18/Z_10 ), .CK(clock), .RN(n1636), 
        .Q(\U3/U1/DATA1_10 ) );
  DFFR_X2 \scratchVal_FS_reg[9]  ( .D(\U18/Z_9 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_9 ) );
  DFFR_X2 \scratchVal_FS_reg[8]  ( .D(\U18/Z_8 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_8 ) );
  DFFR_X2 \scratchVal_FS_reg[7]  ( .D(\U18/Z_7 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_7 ) );
  DFFR_X2 \scratchVal_FS_reg[6]  ( .D(\U18/Z_6 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_6 ) );
  DFFR_X2 \scratchVal_FS_reg[5]  ( .D(\U18/Z_5 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_5 ) );
  DFFR_X2 \scratchVal_FS_reg[4]  ( .D(\U18/Z_4 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_4 ) );
  DFFR_X2 \scratchVal_FS_reg[3]  ( .D(\U18/Z_3 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_3 ) );
  DFFR_X2 \scratchVal_FS_reg[2]  ( .D(\U18/Z_2 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_2 ) );
  DFFR_X2 \scratchVal_FS_reg[1]  ( .D(\U18/Z_1 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_1 ) );
  DFFR_X2 \memoryCounter_reg[2]  ( .D(n1944), .CK(clock), .RN(n1625), .Q(
        \U5/DATA1_2 ), .QN(n1887) );
  DFFR_X2 \memoryCounter_reg[12]  ( .D(n1954), .CK(clock), .RN(n1625), .Q(
        \U5/DATA1_12 ), .QN(n1932) );
  DFFR_X2 \memoryCounter_reg[8]  ( .D(n1950), .CK(clock), .RN(n1625), .Q(
        \U5/DATA1_8 ), .QN(n1913) );
  DFFR_X2 \memoryCounter_reg[10]  ( .D(n1952), .CK(clock), .RN(n1625), .Q(
        \U5/DATA1_10 ), .QN(n1922) );
  DFFR_X2 \memoryCounter_reg[6]  ( .D(n1948), .CK(clock), .RN(n1625), .Q(
        \U5/DATA1_6 ), .QN(n1905) );
  DFFR_X2 \memoryCounter_reg[4]  ( .D(n1946), .CK(clock), .RN(n1625), .Q(
        \U5/DATA1_4 ), .QN(n1896) );
  DFFR_X2 \memoryCounter_reg[1]  ( .D(n1943), .CK(clock), .RN(n1626), .Q(
        \U5/DATA1_1 ) );
  DFFR_X2 \memoryCounter_reg[11]  ( .D(n1953), .CK(clock), .RN(n1626), .Q(
        \U5/DATA1_11 ), .QN(n1878) );
  DFFR_X2 \memoryCounter_reg[9]  ( .D(n1951), .CK(clock), .RN(n1626), .Q(
        \U5/DATA1_9 ), .QN(n1876) );
  DFFR_X2 \memoryCounter_reg[7]  ( .D(n1949), .CK(clock), .RN(n1626), .Q(
        \U5/DATA1_7 ), .QN(n1877) );
  DFFR_X2 \memoryCounter_reg[5]  ( .D(n1947), .CK(clock), .RN(n1626), .Q(
        \U5/DATA1_5 ) );
  DFFR_X2 \memoryCounter_reg[3]  ( .D(n1945), .CK(clock), .RN(n1626), .Q(
        \U5/DATA1_3 ) );
  DFFR_X2 \scratchVal_FS_reg[0]  ( .D(\U18/Z_0 ), .CK(clock), .RN(n1636), .Q(
        \U3/U1/DATA1_0 ) );
  OAI21_X2 U3 ( .B1(n1468), .B2(n212), .A(\U12/Z_0 ), .ZN(\U4/Z_5 ) );
  NOR3_X2 U4 ( .A1(n1787), .A2(n1786), .A3(n1785), .ZN(n1793) );
  NOR2_X2 U6 ( .A1(n1784), .A2(n1783), .ZN(n1795) );
  NAND2_X2 U7 ( .A1(n1424), .A2(n1425), .ZN(\U3/U1/Z_0 ) );
  OAI21_X2 U8 ( .B1(n1467), .B2(n212), .A(\U12/Z_0 ), .ZN(\U4/Z_6 ) );
  OAI21_X2 U9 ( .B1(n1466), .B2(n212), .A(\U12/Z_0 ), .ZN(\U4/Z_4 ) );
  NOR2_X4 U10 ( .A1(\U13/DATA1_5 ), .A2(\U13/DATA1_6 ), .ZN(n1358) );
  NOR2_X4 U11 ( .A1(n157), .A2(n159), .ZN(n1359) );
  AND2_X4 U12 ( .A1(n1462), .A2(n1634), .ZN(n1360) );
  NOR2_X4 U13 ( .A1(n157), .A2(\U13/DATA1_5 ), .ZN(n1361) );
  NOR2_X4 U15 ( .A1(n159), .A2(\U13/DATA1_6 ), .ZN(n1362) );
  AND2_X4 U17 ( .A1(n1883), .A2(n212), .ZN(n1363) );
  AND2_X2 U19 ( .A1(n1794), .A2(n1792), .ZN(n1367) );
  AND2_X4 U21 ( .A1(n1875), .A2(n1634), .ZN(n1368) );
  OR2_X4 U23 ( .A1(\U13/DATA1_3 ), .A2(\U13/DATA1_4 ), .ZN(n1369) );
  AND2_X4 U25 ( .A1(\U13/DATA1_4 ), .A2(\U13/DATA1_3 ), .ZN(n1370) );
  AND2_X4 U27 ( .A1(\U13/DATA1_5 ), .A2(n1370), .ZN(n1371) );
  AND2_X4 U28 ( .A1(\U27/DATA1_9 ), .A2(n1623), .ZN(m2WriteAddr[9]) );
  AND2_X4 U29 ( .A1(\U27/DATA1_10 ), .A2(n1623), .ZN(m2WriteAddr[10]) );
  AND2_X4 U30 ( .A1(\U27/DATA1_11 ), .A2(n1623), .ZN(m2WriteAddr[11]) );
  AND2_X4 U31 ( .A1(\U27/DATA1_13 ), .A2(n1623), .ZN(m2WriteAddr[13]) );
  AND2_X4 U32 ( .A1(\U27/DATA1_15 ), .A2(n1623), .ZN(m2WriteAddr[15]) );
  AND2_X4 U34 ( .A1(\U29/DATA1_8 ), .A2(n1623), .ZN(m2ReadAddr[8]) );
  AND2_X4 U35 ( .A1(n1632), .A2(\U29/DATA1_9 ), .ZN(m2ReadAddr[9]) );
  AND2_X4 U36 ( .A1(\U29/DATA1_10 ), .A2(n1623), .ZN(m2ReadAddr[10]) );
  AND2_X4 U37 ( .A1(\U29/DATA1_12 ), .A2(n1623), .ZN(m2ReadAddr[12]) );
  AND2_X4 U38 ( .A1(\U29/DATA1_14 ), .A2(n1623), .ZN(m2ReadAddr[14]) );
  AND2_X4 U39 ( .A1(\U27/DATA1_8 ), .A2(n1365), .ZN(m2WriteAddr[8]) );
  AND2_X4 U40 ( .A1(\U27/DATA1_12 ), .A2(n1632), .ZN(m2WriteAddr[12]) );
  AND2_X4 U41 ( .A1(\U27/DATA1_14 ), .A2(n1632), .ZN(m2WriteAddr[14]) );
  AND2_X4 U42 ( .A1(\U29/DATA1_11 ), .A2(n1632), .ZN(m2ReadAddr[11]) );
  AND2_X4 U43 ( .A1(\U29/DATA1_13 ), .A2(n1632), .ZN(m2ReadAddr[13]) );
  AND2_X4 U44 ( .A1(\U29/DATA1_15 ), .A2(n1632), .ZN(m2ReadAddr[15]) );
  OAI21_X2 U45 ( .B1(n44), .B2(n1365), .A(n271), .ZN(\U27/Z_5 ) );
  OR2_X1 U54 ( .A1(n1635), .A2(\U14/DATA1_21 ), .ZN(n1399) );
  OR2_X1 U55 ( .A1(n1635), .A2(\U14/DATA1_29 ), .ZN(n1400) );
  OR2_X1 U56 ( .A1(n1635), .A2(\U14/DATA1_23 ), .ZN(n1401) );
  NOR2_X1 U58 ( .A1(\U3/U1/Z_0 ), .A2(n1635), .ZN(n1403) );
  XNOR2_X2 U59 ( .A(n1749), .B(n1742), .ZN(n1743) );
  XNOR2_X2 U60 ( .A(n1404), .B(n1847), .ZN(\U14/DATA1_29 ) );
  XOR2_X2 U61 ( .A(n1862), .B(n1863), .Z(n1416) );
  INV_X4 U62 ( .A(n1421), .ZN(\U14/DATA1_31 ) );
  NAND2_X1 U63 ( .A1(n1449), .A2(n1851), .ZN(n1854) );
  NAND2_X1 U64 ( .A1(n1843), .A2(n1842), .ZN(n1404) );
  OR2_X1 U65 ( .A1(n1786), .A2(n1406), .ZN(n1407) );
  INV_X4 U66 ( .A(n1453), .ZN(n1405) );
  INV_X4 U67 ( .A(n1794), .ZN(n1406) );
  NOR2_X2 U68 ( .A1(n1411), .A2(n1409), .ZN(n1408) );
  INV_X4 U69 ( .A(n1408), .ZN(n1777) );
  OR2_X1 U70 ( .A1(n1406), .A2(n1410), .ZN(n1411) );
  INV_X4 U71 ( .A(n1457), .ZN(n1409) );
  INV_X1 U72 ( .A(n1781), .ZN(n1410) );
  NOR2_X2 U73 ( .A1(n1409), .A2(n1410), .ZN(n1453) );
  NAND2_X2 U74 ( .A1(n1837), .A2(n1830), .ZN(n1414) );
  NAND2_X2 U75 ( .A1(n1412), .A2(n1413), .ZN(n1415) );
  NAND2_X2 U76 ( .A1(n1414), .A2(n1415), .ZN(n1831) );
  INV_X4 U77 ( .A(n1837), .ZN(n1412) );
  INV_X4 U78 ( .A(n1830), .ZN(n1413) );
  NAND3_X2 U79 ( .A1(n1367), .A2(n1795), .A3(n1793), .ZN(n1439) );
  NOR3_X2 U80 ( .A1(n1829), .A2(n1828), .A3(n1827), .ZN(n1830) );
  AND2_X4 U81 ( .A1(n1790), .A2(n1422), .ZN(n1417) );
  AND2_X2 U82 ( .A1(n1460), .A2(n1763), .ZN(n1457) );
  INV_X2 U83 ( .A(n1778), .ZN(n1422) );
  INV_X4 U84 ( .A(n1714), .ZN(n1431) );
  NAND2_X2 U85 ( .A1(n1634), .A2(n1416), .ZN(n1470) );
  NOR2_X2 U86 ( .A1(n1417), .A2(n1418), .ZN(\U14/Z_20 ) );
  NAND2_X1 U87 ( .A1(n1423), .A2(start), .ZN(n1418) );
  INV_X2 U88 ( .A(n1871), .ZN(n1630) );
  INV_X8 U89 ( .A(n1630), .ZN(n1628) );
  NAND2_X1 U90 ( .A1(n1789), .A2(n1778), .ZN(n1423) );
  NOR2_X2 U91 ( .A1(n1405), .A2(n1407), .ZN(n1778) );
  OR2_X2 U92 ( .A1(n1716), .A2(n1715), .ZN(n1446) );
  XNOR2_X1 U93 ( .A(n1747), .B(n1447), .ZN(n1720) );
  NAND2_X4 U94 ( .A1(n1814), .A2(n1819), .ZN(n1827) );
  NAND3_X4 U95 ( .A1(n1753), .A2(n1752), .A3(n1751), .ZN(n1785) );
  NAND2_X1 U96 ( .A1(n1786), .A2(n1777), .ZN(n1419) );
  NAND2_X2 U97 ( .A1(n1773), .A2(n1408), .ZN(n1420) );
  NAND2_X2 U98 ( .A1(n1419), .A2(n1420), .ZN(n1774) );
  OR2_X2 U99 ( .A1(n1617), .A2(n1618), .ZN(n1862) );
  XNOR2_X2 U100 ( .A(n1854), .B(n1852), .ZN(n1421) );
  XNOR2_X1 U101 ( .A(n1781), .B(n1457), .ZN(n1764) );
  AND3_X2 U102 ( .A1(n1464), .A2(n1465), .A3(n1366), .ZN(n1669) );
  NAND3_X2 U103 ( .A1(n1430), .A2(n1781), .A3(n1782), .ZN(n1784) );
  NAND2_X4 U104 ( .A1(n1441), .A2(n1668), .ZN(n1672) );
  NAND2_X1 U105 ( .A1(n1449), .A2(n1851), .ZN(n1617) );
  XNOR2_X1 U106 ( .A(n1851), .B(n1449), .ZN(n1848) );
  INV_X2 U107 ( .A(n1442), .ZN(n1787) );
  NAND2_X2 U108 ( .A1(\U3/U1/DATA1_0 ), .A2(n1630), .ZN(n1424) );
  NAND2_X1 U109 ( .A1(n1673), .A2(n1871), .ZN(n1425) );
  INV_X16 U110 ( .A(n1672), .ZN(n1871) );
  INV_X4 U111 ( .A(\U3/U1/Z_0 ), .ZN(n1432) );
  XNOR2_X1 U112 ( .A(n1713), .B(n1458), .ZN(n1685) );
  AND2_X2 U113 ( .A1(n1458), .A2(n1713), .ZN(n1461) );
  INV_X4 U114 ( .A(n1713), .ZN(n1433) );
  INV_X2 U115 ( .A(n1712), .ZN(n1434) );
  BUF_X4 U116 ( .A(\U5/DATA1_0 ), .Z(m3WriteAddr[0]) );
  BUF_X4 U117 ( .A(\U5/DATA1_1 ), .Z(m3WriteAddr[1]) );
  BUF_X4 U118 ( .A(\U5/DATA1_2 ), .Z(m3WriteAddr[2]) );
  BUF_X4 U119 ( .A(\U5/DATA1_3 ), .Z(m3WriteAddr[3]) );
  BUF_X4 U120 ( .A(\U5/DATA1_4 ), .Z(m3WriteAddr[4]) );
  BUF_X4 U121 ( .A(\U5/DATA1_5 ), .Z(m3WriteAddr[5]) );
  BUF_X4 U122 ( .A(\U5/DATA1_6 ), .Z(m3WriteAddr[6]) );
  BUF_X4 U123 ( .A(\U5/DATA1_7 ), .Z(m3WriteAddr[7]) );
  BUF_X4 U124 ( .A(\U5/DATA1_8 ), .Z(m3WriteAddr[8]) );
  BUF_X4 U125 ( .A(\U5/DATA1_9 ), .Z(m3WriteAddr[9]) );
  BUF_X4 U126 ( .A(\U5/DATA1_10 ), .Z(m3WriteAddr[10]) );
  BUF_X4 U127 ( .A(\U5/DATA1_11 ), .Z(m3WriteAddr[11]) );
  BUF_X4 U128 ( .A(\U5/DATA1_12 ), .Z(m3WriteAddr[12]) );
  BUF_X4 U129 ( .A(\U5/DATA1_13 ), .Z(m3WriteAddr[13]) );
  BUF_X4 U130 ( .A(\U5/DATA1_14 ), .Z(m3WriteAddr[14]) );
  BUF_X4 U131 ( .A(inputBaseOffset), .Z(m3WriteAddr[15]) );
  BUF_X4 U132 ( .A(\U36/DATA2_0 ), .Z(m3WriteBus[0]) );
  BUF_X4 U133 ( .A(\U36/DATA2_1 ), .Z(m3WriteBus[1]) );
  BUF_X4 U134 ( .A(\U36/DATA2_2 ), .Z(m3WriteBus[2]) );
  BUF_X4 U135 ( .A(\U36/DATA2_3 ), .Z(m3WriteBus[3]) );
  BUF_X4 U136 ( .A(\U36/DATA2_4 ), .Z(m3WriteBus[4]) );
  BUF_X4 U137 ( .A(\U36/DATA2_5 ), .Z(m3WriteBus[5]) );
  BUF_X4 U138 ( .A(\U36/DATA2_6 ), .Z(m3WriteBus[6]) );
  BUF_X4 U139 ( .A(\U36/DATA2_7 ), .Z(m3WriteBus[7]) );
  BUF_X4 U140 ( .A(\U36/DATA2_8 ), .Z(m3WriteBus[8]) );
  BUF_X4 U141 ( .A(\U36/DATA2_9 ), .Z(m3WriteBus[9]) );
  BUF_X4 U142 ( .A(\U36/DATA2_10 ), .Z(m3WriteBus[10]) );
  BUF_X4 U143 ( .A(\U36/DATA2_11 ), .Z(m3WriteBus[11]) );
  BUF_X4 U144 ( .A(\U36/DATA2_12 ), .Z(m3WriteBus[12]) );
  BUF_X4 U145 ( .A(\U36/DATA2_13 ), .Z(m3WriteBus[13]) );
  BUF_X4 U146 ( .A(\U36/DATA2_14 ), .Z(m3WriteBus[14]) );
  BUF_X4 U147 ( .A(\U36/DATA2_15 ), .Z(m3WriteBus[15]) );
  BUF_X4 U148 ( .A(\U36/DATA2_16 ), .Z(m3WriteBus[16]) );
  BUF_X4 U149 ( .A(\U36/DATA2_17 ), .Z(m3WriteBus[17]) );
  BUF_X4 U150 ( .A(\U36/DATA2_18 ), .Z(m3WriteBus[18]) );
  BUF_X4 U151 ( .A(\U36/DATA2_19 ), .Z(m3WriteBus[19]) );
  BUF_X4 U152 ( .A(\U36/DATA2_20 ), .Z(m3WriteBus[20]) );
  BUF_X4 U153 ( .A(\U36/DATA2_21 ), .Z(m3WriteBus[21]) );
  BUF_X4 U154 ( .A(\U36/DATA2_22 ), .Z(m3WriteBus[22]) );
  BUF_X4 U155 ( .A(\U36/DATA2_23 ), .Z(m3WriteBus[23]) );
  BUF_X4 U156 ( .A(\U36/DATA2_24 ), .Z(m3WriteBus[24]) );
  BUF_X4 U157 ( .A(\U36/DATA2_25 ), .Z(m3WriteBus[25]) );
  BUF_X4 U158 ( .A(\U36/DATA2_26 ), .Z(m3WriteBus[26]) );
  BUF_X4 U159 ( .A(\U36/DATA2_27 ), .Z(m3WriteBus[27]) );
  BUF_X4 U160 ( .A(\U36/DATA2_28 ), .Z(m3WriteBus[28]) );
  BUF_X4 U161 ( .A(\U36/DATA2_29 ), .Z(m3WriteBus[29]) );
  BUF_X4 U163 ( .A(\U36/DATA2_30 ), .Z(m3WriteBus[30]) );
  BUF_X4 U165 ( .A(\U36/DATA2_31 ), .Z(m3WriteBus[31]) );
  BUF_X4 U167 ( .A(\U36/DATA2_32 ), .Z(m3WriteBus[32]) );
  BUF_X4 U169 ( .A(\U36/DATA2_33 ), .Z(m3WriteBus[33]) );
  BUF_X4 U171 ( .A(\U36/DATA2_34 ), .Z(m3WriteBus[34]) );
  BUF_X4 U173 ( .A(\U36/DATA2_35 ), .Z(m3WriteBus[35]) );
  BUF_X4 U174 ( .A(\U36/DATA2_36 ), .Z(m3WriteBus[36]) );
  BUF_X4 U175 ( .A(\U36/DATA2_37 ), .Z(m3WriteBus[37]) );
  BUF_X4 U176 ( .A(\U36/DATA2_38 ), .Z(m3WriteBus[38]) );
  BUF_X4 U177 ( .A(\U36/DATA2_39 ), .Z(m3WriteBus[39]) );
  BUF_X4 U178 ( .A(\U36/DATA2_40 ), .Z(m3WriteBus[40]) );
  BUF_X4 U179 ( .A(\U36/DATA2_41 ), .Z(m3WriteBus[41]) );
  BUF_X4 U180 ( .A(\U36/DATA2_42 ), .Z(m3WriteBus[42]) );
  BUF_X4 U181 ( .A(\U36/DATA2_43 ), .Z(m3WriteBus[43]) );
  BUF_X4 U182 ( .A(\U36/DATA2_44 ), .Z(m3WriteBus[44]) );
  BUF_X4 U183 ( .A(\U36/DATA2_45 ), .Z(m3WriteBus[45]) );
  BUF_X4 U184 ( .A(\U36/DATA2_46 ), .Z(m3WriteBus[46]) );
  BUF_X4 U185 ( .A(\U36/DATA2_47 ), .Z(m3WriteBus[47]) );
  BUF_X4 U187 ( .A(\U36/DATA2_48 ), .Z(m3WriteBus[48]) );
  BUF_X4 U189 ( .A(\U36/DATA2_49 ), .Z(m3WriteBus[49]) );
  BUF_X4 U191 ( .A(\U36/DATA2_50 ), .Z(m3WriteBus[50]) );
  BUF_X4 U192 ( .A(\U36/DATA2_51 ), .Z(m3WriteBus[51]) );
  BUF_X4 U193 ( .A(\U36/DATA2_52 ), .Z(m3WriteBus[52]) );
  BUF_X4 U194 ( .A(\U36/DATA2_53 ), .Z(m3WriteBus[53]) );
  BUF_X4 U195 ( .A(\U36/DATA2_54 ), .Z(m3WriteBus[54]) );
  BUF_X4 U197 ( .A(\U36/DATA2_55 ), .Z(m3WriteBus[55]) );
  BUF_X4 U199 ( .A(\U36/DATA2_56 ), .Z(m3WriteBus[56]) );
  BUF_X4 U201 ( .A(\U36/DATA2_57 ), .Z(m3WriteBus[57]) );
  BUF_X4 U203 ( .A(\U36/DATA2_58 ), .Z(m3WriteBus[58]) );
  BUF_X4 U205 ( .A(\U36/DATA2_59 ), .Z(m3WriteBus[59]) );
  BUF_X4 U207 ( .A(\U36/DATA2_60 ), .Z(m3WriteBus[60]) );
  BUF_X4 U208 ( .A(\U36/DATA2_61 ), .Z(m3WriteBus[61]) );
  BUF_X4 U209 ( .A(\U36/DATA2_62 ), .Z(m3WriteBus[62]) );
  BUF_X4 U210 ( .A(\U36/DATA2_63 ), .Z(m3WriteBus[63]) );
  BUF_X4 U211 ( .A(\U36/DATA2_64 ), .Z(m3WriteBus[64]) );
  BUF_X4 U212 ( .A(\U36/DATA2_65 ), .Z(m3WriteBus[65]) );
  BUF_X4 U213 ( .A(\U36/DATA2_66 ), .Z(m3WriteBus[66]) );
  BUF_X4 U214 ( .A(\U36/DATA2_67 ), .Z(m3WriteBus[67]) );
  BUF_X4 U215 ( .A(\U36/DATA2_68 ), .Z(m3WriteBus[68]) );
  BUF_X4 U216 ( .A(\U36/DATA2_69 ), .Z(m3WriteBus[69]) );
  BUF_X4 U217 ( .A(\U36/DATA2_70 ), .Z(m3WriteBus[70]) );
  BUF_X4 U218 ( .A(\U36/DATA1_7 ), .Z(m3WriteBus[71]) );
  BUF_X4 U219 ( .A(\U36/DATA1_8 ), .Z(m3WriteBus[72]) );
  BUF_X4 U221 ( .A(\U36/DATA1_9 ), .Z(m3WriteBus[73]) );
  BUF_X4 U223 ( .A(\U36/DATA1_10 ), .Z(m3WriteBus[74]) );
  BUF_X4 U225 ( .A(\U36/DATA1_11 ), .Z(m3WriteBus[75]) );
  BUF_X4 U227 ( .A(\U36/DATA1_12 ), .Z(m3WriteBus[76]) );
  BUF_X4 U229 ( .A(\U36/DATA1_13 ), .Z(m3WriteBus[77]) );
  BUF_X4 U231 ( .A(\U36/DATA1_14 ), .Z(m3WriteBus[78]) );
  BUF_X4 U233 ( .A(\U36/DATA1_15 ), .Z(m3WriteBus[79]) );
  BUF_X4 U235 ( .A(\U36/DATA1_16 ), .Z(m3WriteBus[80]) );
  BUF_X4 U237 ( .A(\U36/DATA1_17 ), .Z(m3WriteBus[81]) );
  BUF_X4 U239 ( .A(\U36/DATA1_18 ), .Z(m3WriteBus[82]) );
  BUF_X4 U241 ( .A(\U36/DATA1_19 ), .Z(m3WriteBus[83]) );
  BUF_X4 U243 ( .A(\U36/DATA1_20 ), .Z(m3WriteBus[84]) );
  BUF_X4 U245 ( .A(\U36/DATA1_21 ), .Z(m3WriteBus[85]) );
  BUF_X4 U247 ( .A(\U36/DATA1_22 ), .Z(m3WriteBus[86]) );
  BUF_X4 U249 ( .A(\U36/DATA1_23 ), .Z(m3WriteBus[87]) );
  BUF_X4 U251 ( .A(\U36/DATA1_24 ), .Z(m3WriteBus[88]) );
  BUF_X4 U253 ( .A(\U36/DATA1_25 ), .Z(m3WriteBus[89]) );
  BUF_X4 U255 ( .A(\U36/DATA1_26 ), .Z(m3WriteBus[90]) );
  BUF_X4 U257 ( .A(\U36/DATA1_27 ), .Z(m3WriteBus[91]) );
  BUF_X4 U259 ( .A(\U36/DATA1_28 ), .Z(m3WriteBus[92]) );
  BUF_X4 U261 ( .A(\U36/DATA1_29 ), .Z(m3WriteBus[93]) );
  BUF_X4 U263 ( .A(\U36/DATA1_30 ), .Z(m3WriteBus[94]) );
  BUF_X4 U265 ( .A(\U36/DATA1_31 ), .Z(m3WriteBus[95]) );
  BUF_X4 U267 ( .A(\U36/DATA1_32 ), .Z(m3WriteBus[96]) );
  BUF_X4 U269 ( .A(\U36/DATA1_33 ), .Z(m3WriteBus[97]) );
  BUF_X4 U271 ( .A(\U36/DATA1_34 ), .Z(m3WriteBus[98]) );
  BUF_X4 U273 ( .A(\U36/DATA1_35 ), .Z(m3WriteBus[99]) );
  BUF_X4 U275 ( .A(\U36/DATA1_36 ), .Z(m3WriteBus[100]) );
  BUF_X4 U277 ( .A(\U36/DATA1_37 ), .Z(m3WriteBus[101]) );
  BUF_X4 U279 ( .A(\U36/DATA1_38 ), .Z(m3WriteBus[102]) );
  BUF_X4 U281 ( .A(\U36/DATA1_39 ), .Z(m3WriteBus[103]) );
  BUF_X4 U283 ( .A(\U36/DATA1_40 ), .Z(m3WriteBus[104]) );
  BUF_X4 U285 ( .A(\U36/DATA1_41 ), .Z(m3WriteBus[105]) );
  BUF_X4 U287 ( .A(\U36/DATA1_42 ), .Z(m3WriteBus[106]) );
  BUF_X4 U289 ( .A(\U36/DATA1_43 ), .Z(m3WriteBus[107]) );
  BUF_X4 U291 ( .A(\U36/DATA1_44 ), .Z(m3WriteBus[108]) );
  BUF_X4 U293 ( .A(\U36/DATA1_45 ), .Z(m3WriteBus[109]) );
  BUF_X4 U295 ( .A(\U36/DATA1_46 ), .Z(m3WriteBus[110]) );
  BUF_X4 U296 ( .A(\U36/DATA1_47 ), .Z(m3WriteBus[111]) );
  BUF_X4 U297 ( .A(\U36/DATA1_48 ), .Z(m3WriteBus[112]) );
  BUF_X4 U298 ( .A(\U36/DATA1_49 ), .Z(m3WriteBus[113]) );
  BUF_X4 U299 ( .A(\U36/DATA1_50 ), .Z(m3WriteBus[114]) );
  BUF_X4 U300 ( .A(\U36/DATA1_51 ), .Z(m3WriteBus[115]) );
  BUF_X4 U301 ( .A(\U36/DATA1_52 ), .Z(m3WriteBus[116]) );
  BUF_X4 U302 ( .A(\U36/DATA1_53 ), .Z(m3WriteBus[117]) );
  BUF_X4 U303 ( .A(\U36/DATA1_54 ), .Z(m3WriteBus[118]) );
  BUF_X4 U304 ( .A(\U36/DATA1_55 ), .Z(m3WriteBus[119]) );
  BUF_X4 U305 ( .A(\U36/DATA1_56 ), .Z(m3WriteBus[120]) );
  BUF_X4 U306 ( .A(\U36/DATA1_57 ), .Z(m3WriteBus[121]) );
  BUF_X4 U307 ( .A(\U36/DATA1_58 ), .Z(m3WriteBus[122]) );
  BUF_X4 U308 ( .A(\U36/DATA1_59 ), .Z(m3WriteBus[123]) );
  BUF_X4 U309 ( .A(\U36/DATA1_60 ), .Z(m3WriteBus[124]) );
  BUF_X4 U310 ( .A(\U36/DATA1_61 ), .Z(m3WriteBus[125]) );
  BUF_X4 U311 ( .A(\U36/DATA1_62 ), .Z(m3WriteBus[126]) );
  BUF_X4 U312 ( .A(\U36/DATA1_63 ), .Z(m3WriteBus[127]) );
  NAND2_X2 U313 ( .A1(n1873), .A2(n1427), .ZN(n1428) );
  NAND2_X2 U314 ( .A1(n1426), .A2(n1872), .ZN(n1429) );
  NAND2_X2 U315 ( .A1(n1428), .A2(n1429), .ZN(n1874) );
  INV_X2 U316 ( .A(n1873), .ZN(n1426) );
  INV_X1 U317 ( .A(n1872), .ZN(n1427) );
  NOR4_X2 U318 ( .A1(n1431), .A2(n1432), .A3(n1433), .A4(n1434), .ZN(n1430) );
  AND4_X2 U319 ( .A1(n1435), .A2(n1436), .A3(n1437), .A4(n1438), .ZN(n1668) );
  XNOR2_X2 U320 ( .A(\U27/DATA2_0 ), .B(\U15/DATA1_0 ), .ZN(n1435) );
  XOR2_X2 U321 ( .A(n48), .B(\U15/DATA1_1 ), .Z(n1436) );
  XNOR2_X2 U322 ( .A(n1666), .B(n47), .ZN(n1437) );
  XNOR2_X2 U324 ( .A(n1667), .B(n46), .ZN(n1438) );
  NAND4_X1 U326 ( .A1(n1795), .A2(n1793), .A3(n1794), .A4(n1792), .ZN(n1798)
         );
  NAND3_X2 U327 ( .A1(n1671), .A2(n1670), .A3(n1669), .ZN(n1440) );
  INV_X4 U330 ( .A(n1440), .ZN(n1441) );
  AND2_X4 U332 ( .A1(n1447), .A2(n1747), .ZN(n1456) );
  AND2_X2 U333 ( .A1(n1448), .A2(n1788), .ZN(n1460) );
  AND2_X4 U336 ( .A1(\U26/DATA1_36 ), .A2(n1623), .ZN(\U26/Z_36 ) );
  AND2_X4 U338 ( .A1(\U26/DATA1_37 ), .A2(n1632), .ZN(\U26/Z_37 ) );
  AND2_X4 U340 ( .A1(\U26/DATA1_38 ), .A2(n1623), .ZN(\U26/Z_38 ) );
  AND2_X4 U341 ( .A1(\U26/DATA1_39 ), .A2(n1632), .ZN(\U26/Z_39 ) );
  AND2_X4 U343 ( .A1(\U26/DATA1_40 ), .A2(n1623), .ZN(\U26/Z_40 ) );
  AND2_X4 U344 ( .A1(\U26/DATA1_41 ), .A2(n1632), .ZN(\U26/Z_41 ) );
  AND2_X4 U345 ( .A1(\U26/DATA1_42 ), .A2(n1623), .ZN(\U26/Z_42 ) );
  AND2_X4 U347 ( .A1(\U26/DATA1_43 ), .A2(n1632), .ZN(\U26/Z_43 ) );
  AND2_X4 U348 ( .A1(\U26/DATA1_44 ), .A2(n1623), .ZN(\U26/Z_44 ) );
  AND2_X4 U349 ( .A1(\U26/DATA1_45 ), .A2(n1632), .ZN(\U26/Z_45 ) );
  AND2_X4 U352 ( .A1(\U26/DATA1_46 ), .A2(n1623), .ZN(\U26/Z_46 ) );
  AND2_X4 U354 ( .A1(\U26/DATA1_47 ), .A2(n1632), .ZN(\U26/Z_47 ) );
  AND2_X4 U355 ( .A1(\U26/DATA1_48 ), .A2(n1623), .ZN(\U26/Z_48 ) );
  AND2_X4 U358 ( .A1(\U26/DATA1_49 ), .A2(n1632), .ZN(\U26/Z_49 ) );
  AND2_X4 U360 ( .A1(\U26/DATA1_50 ), .A2(n1623), .ZN(\U26/Z_50 ) );
  AND2_X4 U362 ( .A1(\U26/DATA1_51 ), .A2(n1632), .ZN(\U26/Z_51 ) );
  AND2_X4 U363 ( .A1(\U26/DATA1_52 ), .A2(n1623), .ZN(\U26/Z_52 ) );
  AND2_X4 U365 ( .A1(\U26/DATA1_53 ), .A2(n1623), .ZN(\U26/Z_53 ) );
  AND2_X4 U366 ( .A1(\U26/DATA1_54 ), .A2(n1632), .ZN(\U26/Z_54 ) );
  AND2_X4 U367 ( .A1(\U26/DATA1_55 ), .A2(n1623), .ZN(\U26/Z_55 ) );
  AND2_X4 U368 ( .A1(\U26/DATA1_56 ), .A2(n1632), .ZN(\U26/Z_56 ) );
  AND2_X4 U371 ( .A1(\U26/DATA1_57 ), .A2(n1623), .ZN(\U26/Z_57 ) );
  AND2_X4 U373 ( .A1(\U26/DATA1_58 ), .A2(n1632), .ZN(\U26/Z_58 ) );
  AND2_X4 U374 ( .A1(\U26/DATA1_59 ), .A2(n1623), .ZN(\U26/Z_59 ) );
  AND2_X4 U375 ( .A1(\U26/DATA1_60 ), .A2(n1632), .ZN(\U26/Z_60 ) );
  AND2_X4 U377 ( .A1(\U26/DATA1_61 ), .A2(n1623), .ZN(\U26/Z_61 ) );
  AND2_X4 U378 ( .A1(\U26/DATA1_62 ), .A2(n1632), .ZN(\U26/Z_62 ) );
  AND2_X4 U381 ( .A1(\U26/DATA1_63 ), .A2(n1623), .ZN(\U26/Z_63 ) );
  AND2_X4 U383 ( .A1(\U26/DATA1_64 ), .A2(n1632), .ZN(\U26/Z_64 ) );
  AND2_X4 U384 ( .A1(\U26/DATA1_65 ), .A2(n1623), .ZN(\U26/Z_65 ) );
  AND2_X4 U385 ( .A1(\U26/DATA1_66 ), .A2(n1632), .ZN(\U26/Z_66 ) );
  AND2_X4 U387 ( .A1(\U26/DATA1_67 ), .A2(n1623), .ZN(\U26/Z_67 ) );
  AND2_X4 U388 ( .A1(\U26/DATA1_68 ), .A2(n1632), .ZN(\U26/Z_68 ) );
  AND2_X4 U389 ( .A1(\U26/DATA1_69 ), .A2(n1623), .ZN(\U26/Z_69 ) );
  AND2_X4 U391 ( .A1(\U26/DATA1_70 ), .A2(n1632), .ZN(\U26/Z_70 ) );
  AND2_X4 U392 ( .A1(\U26/DATA1_71 ), .A2(n1623), .ZN(\U26/Z_71 ) );
  AND2_X4 U394 ( .A1(\U26/DATA1_72 ), .A2(n1632), .ZN(\U26/Z_72 ) );
  AND2_X4 U395 ( .A1(\U26/DATA1_73 ), .A2(n1623), .ZN(\U26/Z_73 ) );
  AND2_X4 U399 ( .A1(\U26/DATA1_74 ), .A2(n1632), .ZN(\U26/Z_74 ) );
  AND2_X4 U401 ( .A1(\U26/DATA1_75 ), .A2(n1623), .ZN(\U26/Z_75 ) );
  AND2_X4 U402 ( .A1(\U26/DATA1_76 ), .A2(n1632), .ZN(\U26/Z_76 ) );
  AND2_X4 U403 ( .A1(\U26/DATA1_77 ), .A2(n1623), .ZN(\U26/Z_77 ) );
  AND2_X4 U404 ( .A1(\U26/DATA1_78 ), .A2(n1632), .ZN(\U26/Z_78 ) );
  AND2_X4 U405 ( .A1(\U26/DATA1_79 ), .A2(n1623), .ZN(\U26/Z_79 ) );
  AND2_X4 U406 ( .A1(\U26/DATA1_80 ), .A2(n1632), .ZN(\U26/Z_80 ) );
  AND2_X4 U407 ( .A1(\U26/DATA1_81 ), .A2(n1623), .ZN(\U26/Z_81 ) );
  AND2_X4 U408 ( .A1(\U26/DATA1_82 ), .A2(n1632), .ZN(\U26/Z_82 ) );
  AND2_X4 U409 ( .A1(\U26/DATA1_83 ), .A2(n1623), .ZN(\U26/Z_83 ) );
  AND2_X4 U410 ( .A1(\U26/DATA1_84 ), .A2(n1632), .ZN(\U26/Z_84 ) );
  AND2_X4 U411 ( .A1(\U26/DATA1_85 ), .A2(n1623), .ZN(\U26/Z_85 ) );
  AND2_X4 U412 ( .A1(\U26/DATA1_86 ), .A2(n1632), .ZN(\U26/Z_86 ) );
  AND2_X4 U413 ( .A1(\U26/DATA1_87 ), .A2(n1623), .ZN(\U26/Z_87 ) );
  AND2_X4 U414 ( .A1(\U26/DATA1_88 ), .A2(n1632), .ZN(\U26/Z_88 ) );
  AND2_X4 U415 ( .A1(\U26/DATA1_89 ), .A2(n1623), .ZN(\U26/Z_89 ) );
  AND2_X4 U416 ( .A1(\U26/DATA1_90 ), .A2(n1632), .ZN(\U26/Z_90 ) );
  AND2_X4 U417 ( .A1(\U26/DATA1_91 ), .A2(n1623), .ZN(\U26/Z_91 ) );
  AND2_X4 U418 ( .A1(\U26/DATA1_92 ), .A2(n1632), .ZN(\U26/Z_92 ) );
  AND2_X4 U419 ( .A1(\U26/DATA1_93 ), .A2(n1623), .ZN(\U26/Z_93 ) );
  AND2_X4 U420 ( .A1(\U26/DATA1_94 ), .A2(n1632), .ZN(\U26/Z_94 ) );
  AND2_X4 U421 ( .A1(\U26/DATA1_95 ), .A2(n1623), .ZN(\U26/Z_95 ) );
  AND2_X4 U422 ( .A1(\U26/DATA1_96 ), .A2(n1632), .ZN(\U26/Z_96 ) );
  AND2_X4 U423 ( .A1(\U26/DATA1_97 ), .A2(n1623), .ZN(\U26/Z_97 ) );
  AND2_X4 U424 ( .A1(\U26/DATA1_98 ), .A2(n1623), .ZN(\U26/Z_98 ) );
  AND2_X4 U425 ( .A1(\U26/DATA1_99 ), .A2(n1632), .ZN(\U26/Z_99 ) );
  AND2_X4 U426 ( .A1(\U26/DATA1_100 ), .A2(n1623), .ZN(\U26/Z_100 ) );
  AND2_X4 U427 ( .A1(\U26/DATA1_101 ), .A2(n1623), .ZN(\U26/Z_101 ) );
  AND2_X4 U428 ( .A1(\U26/DATA1_102 ), .A2(n1632), .ZN(\U26/Z_102 ) );
  AND2_X4 U429 ( .A1(\U26/DATA1_103 ), .A2(n1623), .ZN(\U26/Z_103 ) );
  AND2_X4 U430 ( .A1(\U26/DATA1_104 ), .A2(n1632), .ZN(\U26/Z_104 ) );
  AND2_X4 U431 ( .A1(\U26/DATA1_105 ), .A2(n1623), .ZN(\U26/Z_105 ) );
  AND2_X4 U432 ( .A1(\U26/DATA1_106 ), .A2(n1632), .ZN(\U26/Z_106 ) );
  AND2_X4 U433 ( .A1(\U26/DATA1_107 ), .A2(n1623), .ZN(\U26/Z_107 ) );
  AND2_X4 U434 ( .A1(\U26/DATA1_108 ), .A2(n1632), .ZN(\U26/Z_108 ) );
  AND2_X4 U435 ( .A1(\U26/DATA1_109 ), .A2(n1632), .ZN(\U26/Z_109 ) );
  AND2_X4 U436 ( .A1(\U26/DATA1_110 ), .A2(n1623), .ZN(\U26/Z_110 ) );
  AND2_X4 U437 ( .A1(\U26/DATA1_111 ), .A2(n1632), .ZN(\U26/Z_111 ) );
  AND2_X4 U438 ( .A1(\U26/DATA1_112 ), .A2(n1623), .ZN(\U26/Z_112 ) );
  AND2_X4 U439 ( .A1(\U26/DATA1_113 ), .A2(n1632), .ZN(\U26/Z_113 ) );
  AND2_X4 U440 ( .A1(\U26/DATA1_114 ), .A2(n1623), .ZN(\U26/Z_114 ) );
  AND2_X4 U441 ( .A1(\U26/DATA1_115 ), .A2(n1632), .ZN(\U26/Z_115 ) );
  AND2_X4 U442 ( .A1(\U26/DATA1_116 ), .A2(n1623), .ZN(\U26/Z_116 ) );
  AND2_X4 U443 ( .A1(\U26/DATA1_117 ), .A2(n1632), .ZN(\U26/Z_117 ) );
  AND2_X4 U444 ( .A1(\U26/DATA1_118 ), .A2(n1623), .ZN(\U26/Z_118 ) );
  AND2_X4 U445 ( .A1(\U26/DATA1_119 ), .A2(n1632), .ZN(\U26/Z_119 ) );
  AND2_X4 U446 ( .A1(\U26/DATA1_120 ), .A2(n1623), .ZN(\U26/Z_120 ) );
  AND2_X4 U447 ( .A1(\U26/DATA1_121 ), .A2(n1632), .ZN(\U26/Z_121 ) );
  AND2_X4 U448 ( .A1(\U26/DATA1_122 ), .A2(n1623), .ZN(\U26/Z_122 ) );
  AND2_X4 U449 ( .A1(\U26/DATA1_123 ), .A2(n1632), .ZN(\U26/Z_123 ) );
  AND2_X4 U450 ( .A1(\U26/DATA1_124 ), .A2(n1623), .ZN(\U26/Z_124 ) );
  AND2_X4 U451 ( .A1(\U26/DATA1_125 ), .A2(n1632), .ZN(\U26/Z_125 ) );
  AND2_X4 U452 ( .A1(\U26/DATA1_126 ), .A2(n1623), .ZN(\U26/Z_126 ) );
  AND2_X4 U453 ( .A1(\U26/DATA1_127 ), .A2(n1632), .ZN(\U26/Z_127 ) );
  XNOR2_X1 U454 ( .A(n1620), .B(n1838), .ZN(\U14/DATA1_23 ) );
  AND2_X2 U455 ( .A1(n1430), .A2(n1442), .ZN(n1447) );
  INV_X4 U463 ( .A(n1847), .ZN(n1450) );
  AND2_X4 U464 ( .A1(n1712), .A2(\U3/U1/Z_0 ), .ZN(n1451) );
  XOR2_X1 U465 ( .A(n1834), .B(n1800), .Z(n1801) );
  XNOR2_X1 U466 ( .A(n1813), .B(n1819), .ZN(\U14/DATA1_25 ) );
  INV_X4 U467 ( .A(n1719), .ZN(n1443) );
  INV_X4 U468 ( .A(n1718), .ZN(n1444) );
  INV_X4 U469 ( .A(n1717), .ZN(n1445) );
  INV_X2 U470 ( .A(n400), .ZN(n1965) );
  INV_X2 U471 ( .A(n382), .ZN(n1970) );
  NOR4_X2 U472 ( .A1(n1446), .A2(n1443), .A3(n1444), .A4(n1445), .ZN(n1442) );
  INV_X4 U473 ( .A(n1360), .ZN(n1627) );
  INV_X8 U474 ( .A(n1631), .ZN(n1623) );
  INV_X16 U475 ( .A(n1637), .ZN(n1636) );
  INV_X4 U476 ( .A(n1637), .ZN(n1625) );
  INV_X4 U477 ( .A(n1637), .ZN(n1624) );
  INV_X4 U478 ( .A(n1637), .ZN(n1626) );
  INV_X4 U479 ( .A(n1630), .ZN(n1629) );
  AND3_X2 U480 ( .A1(n1782), .A2(n1754), .A3(n1447), .ZN(n1448) );
  INV_X4 U481 ( .A(rst_n), .ZN(n1637) );
  NAND2_X2 U482 ( .A1(n1368), .A2(n211), .ZN(n209) );
  INV_X1 U483 ( .A(n1834), .ZN(n1621) );
  NOR2_X1 U484 ( .A1(n1854), .A2(n1852), .ZN(n1622) );
  NAND2_X2 U485 ( .A1(n1620), .A2(n1806), .ZN(n1824) );
  XNOR2_X2 U486 ( .A(n1717), .B(n1707), .ZN(n1708) );
  NOR2_X2 U487 ( .A1(n1846), .A2(n1450), .ZN(n1449) );
  AND2_X1 U488 ( .A1(n1456), .A2(n1751), .ZN(n1452) );
  AND2_X1 U489 ( .A1(n1452), .A2(n1752), .ZN(n1454) );
  AND2_X1 U490 ( .A1(n1459), .A2(n1714), .ZN(n1455) );
  AND2_X1 U491 ( .A1(n1451), .A2(n1684), .ZN(n1458) );
  AND2_X1 U492 ( .A1(n1461), .A2(n1693), .ZN(n1459) );
  AND3_X2 U493 ( .A1(n1661), .A2(n1660), .A3(n1659), .ZN(n1462) );
  INV_X4 U494 ( .A(n1635), .ZN(n1634) );
  INV_X4 U495 ( .A(n1632), .ZN(n1631) );
  NAND4_X2 U496 ( .A1(n455), .A2(n456), .A3(n453), .A4(n454), .ZN(n1772) );
  AOI22_X2 U497 ( .A1(\U36/DATA1_44 ), .A2(n1359), .B1(\U36/DATA2_12 ), .B2(
        n1358), .ZN(n400) );
  AOI22_X2 U498 ( .A1(\U36/DATA1_46 ), .A2(n1359), .B1(\U36/DATA2_14 ), .B2(
        n1358), .ZN(n382) );
  AOI22_X2 U499 ( .A1(\U36/DATA1_42 ), .A2(n1359), .B1(\U36/DATA2_10 ), .B2(
        n1358), .ZN(n378) );
  AOI22_X2 U500 ( .A1(\U36/DATA1_43 ), .A2(n1359), .B1(\U36/DATA2_11 ), .B2(
        n1358), .ZN(n433) );
  AOI22_X2 U501 ( .A1(\U36/DATA1_60 ), .A2(n1359), .B1(\U36/DATA2_28 ), .B2(
        n1358), .ZN(n401) );
  AOI22_X2 U502 ( .A1(\U36/DATA1_62 ), .A2(n1359), .B1(\U36/DATA2_30 ), .B2(
        n1358), .ZN(n383) );
  AOI22_X2 U503 ( .A1(\U36/DATA1_58 ), .A2(n1359), .B1(\U36/DATA2_26 ), .B2(
        n1358), .ZN(n379) );
  AOI22_X2 U504 ( .A1(\U36/DATA1_59 ), .A2(n1359), .B1(\U36/DATA2_27 ), .B2(
        n1358), .ZN(n434) );
  AOI22_X2 U505 ( .A1(n1361), .A2(\U36/DATA2_68 ), .B1(n1362), .B2(
        \U36/DATA2_36 ), .ZN(n405) );
  AOI22_X2 U506 ( .A1(\U36/DATA1_34 ), .A2(n1359), .B1(\U36/DATA2_2 ), .B2(
        n1358), .ZN(n372) );
  AOI22_X2 U507 ( .A1(\U36/DATA1_35 ), .A2(n1359), .B1(\U36/DATA2_3 ), .B2(
        n1358), .ZN(n428) );
  AOI22_X2 U508 ( .A1(\U36/DATA2_55 ), .A2(n1362), .B1(\U36/DATA1_23 ), .B2(
        n1361), .ZN(n447) );
  AOI22_X2 U509 ( .A1(\U36/DATA1_55 ), .A2(n1359), .B1(\U36/DATA2_23 ), .B2(
        n1358), .ZN(n448) );
  OR2_X1 U510 ( .A1(n1463), .A2(n1937), .ZN(n1939) );
  AOI22_X2 U511 ( .A1(\U36/DATA2_50 ), .A2(n1362), .B1(\U36/DATA1_18 ), .B2(
        n1361), .ZN(n374) );
  AOI22_X2 U512 ( .A1(\U36/DATA2_51 ), .A2(n1362), .B1(\U36/DATA1_19 ), .B2(
        n1361), .ZN(n429) );
  AOI22_X2 U514 ( .A1(\U36/DATA2_52 ), .A2(n1362), .B1(\U36/DATA1_20 ), .B2(
        n1361), .ZN(n402) );
  AOI22_X2 U515 ( .A1(\U36/DATA2_54 ), .A2(n1362), .B1(\U36/DATA1_22 ), .B2(
        n1361), .ZN(n384) );
  AOI22_X2 U516 ( .A1(\U36/DATA1_51 ), .A2(n1359), .B1(\U36/DATA2_19 ), .B2(
        n1358), .ZN(n430) );
  AOI22_X2 U517 ( .A1(\U36/DATA1_50 ), .A2(n1359), .B1(\U36/DATA2_18 ), .B2(
        n1358), .ZN(n375) );
  AOI22_X2 U518 ( .A1(\U36/DATA1_52 ), .A2(n1359), .B1(\U36/DATA2_20 ), .B2(
        n1358), .ZN(n403) );
  AOI22_X2 U519 ( .A1(\U36/DATA1_54 ), .A2(n1359), .B1(\U36/DATA2_22 ), .B2(
        n1358), .ZN(n385) );
  AOI22_X2 U520 ( .A1(\U36/DATA1_48 ), .A2(n1359), .B1(\U36/DATA2_16 ), .B2(
        n1358), .ZN(n392) );
  AOI22_X2 U521 ( .A1(\U36/DATA1_49 ), .A2(n1359), .B1(\U36/DATA2_17 ), .B2(
        n1358), .ZN(n424) );
  AOI22_X2 U522 ( .A1(\U36/DATA1_53 ), .A2(n1359), .B1(\U36/DATA2_21 ), .B2(
        n1358), .ZN(n415) );
  AOI22_X2 U524 ( .A1(\U36/DATA2_48 ), .A2(n1362), .B1(\U36/DATA1_16 ), .B2(
        n1361), .ZN(n391) );
  AOI22_X2 U525 ( .A1(\U36/DATA2_49 ), .A2(n1362), .B1(\U36/DATA1_17 ), .B2(
        n1361), .ZN(n423) );
  AOI22_X2 U526 ( .A1(\U36/DATA2_53 ), .A2(n1362), .B1(\U36/DATA1_21 ), .B2(
        n1361), .ZN(n414) );
  AOI21_X2 U527 ( .B1(n441), .B2(n442), .A(\U13/DATA1_3 ), .ZN(n437) );
  AOI22_X2 U528 ( .A1(\U36/DATA2_39 ), .A2(n1362), .B1(\U36/DATA1_7 ), .B2(
        n1361), .ZN(n441) );
  AOI22_X2 U529 ( .A1(\U36/DATA1_39 ), .A2(n1359), .B1(\U36/DATA2_7 ), .B2(
        n1358), .ZN(n442) );
  AOI21_X2 U530 ( .B1(n439), .B2(n440), .A(n167), .ZN(n438) );
  AOI22_X2 U531 ( .A1(\U36/DATA2_47 ), .A2(n1362), .B1(\U36/DATA1_15 ), .B2(
        n1361), .ZN(n439) );
  AOI22_X2 U532 ( .A1(\U36/DATA1_47 ), .A2(n1359), .B1(\U36/DATA2_15 ), .B2(
        n1358), .ZN(n440) );
  AOI21_X2 U533 ( .B1(n445), .B2(n446), .A(n167), .ZN(n444) );
  AOI22_X2 U534 ( .A1(\U36/DATA2_63 ), .A2(n1362), .B1(\U36/DATA1_31 ), .B2(
        n1361), .ZN(n445) );
  AOI22_X2 U535 ( .A1(\U36/DATA1_63 ), .A2(n1359), .B1(\U36/DATA2_31 ), .B2(
        n1358), .ZN(n446) );
  XNOR2_X2 U536 ( .A(n1663), .B(n44), .ZN(n1464) );
  XNOR2_X2 U537 ( .A(n1664), .B(n45), .ZN(n1465) );
  OAI21_X2 U538 ( .B1(n172), .B2(n1363), .A(n1942), .ZN(n511) );
  XOR2_X2 U539 ( .A(n165), .B(\U13/DATA1_3 ), .Z(n1466) );
  OAI21_X2 U540 ( .B1(\U13/DATA1_3 ), .B2(n212), .A(\U12/Z_0 ), .ZN(\U4/Z_3 )
         );
  XOR2_X2 U541 ( .A(n157), .B(n1371), .Z(n1467) );
  XOR2_X2 U542 ( .A(n159), .B(n1370), .Z(n1468) );
  OAI21_X2 U543 ( .B1(n443), .B2(n444), .A(\U13/DATA1_4 ), .ZN(n435) );
  OAI21_X2 U544 ( .B1(n437), .B2(n438), .A(n165), .ZN(n436) );
  AOI21_X2 U545 ( .B1(n447), .B2(n448), .A(\U13/DATA1_3 ), .ZN(n443) );
  AOI22_X2 U546 ( .A1(\U36/DATA2_70 ), .A2(n1361), .B1(\U36/DATA2_38 ), .B2(
        n1362), .ZN(n387) );
  AOI22_X2 U547 ( .A1(\U36/DATA1_40 ), .A2(n1359), .B1(\U36/DATA2_8 ), .B2(
        n1358), .ZN(n396) );
  AOI22_X2 U548 ( .A1(\U36/DATA1_56 ), .A2(n1359), .B1(\U36/DATA2_24 ), .B2(
        n1358), .ZN(n397) );
  AOI22_X2 U549 ( .A1(\U36/DATA1_41 ), .A2(n1359), .B1(\U36/DATA2_9 ), .B2(
        n1358), .ZN(n421) );
  AOI22_X2 U550 ( .A1(\U36/DATA1_57 ), .A2(n1359), .B1(\U36/DATA2_25 ), .B2(
        n1358), .ZN(n422) );
  AOI22_X2 U551 ( .A1(\U36/DATA1_45 ), .A2(n1359), .B1(\U36/DATA2_13 ), .B2(
        n1358), .ZN(n412) );
  AOI22_X2 U552 ( .A1(\U36/DATA1_61 ), .A2(n1359), .B1(\U36/DATA2_29 ), .B2(
        n1358), .ZN(n413) );
  AOI22_X2 U553 ( .A1(\U36/DATA1_32 ), .A2(n1359), .B1(\U36/DATA2_0 ), .B2(
        n1358), .ZN(n390) );
  AOI22_X2 U554 ( .A1(n1361), .A2(\U36/DATA2_65 ), .B1(n1362), .B2(
        \U36/DATA2_33 ), .ZN(n425) );
  AOI22_X2 U555 ( .A1(n1361), .A2(\U36/DATA2_69 ), .B1(n1362), .B2(
        \U36/DATA2_37 ), .ZN(n416) );
  INV_X4 U556 ( .A(start), .ZN(n1635) );
  INV_X4 U557 ( .A(n1633), .ZN(n1632) );
  OAI21_X2 U558 ( .B1(n47), .B2(n1623), .A(n274), .ZN(\U27/Z_2 ) );
  OAI21_X2 U559 ( .B1(n45), .B2(n1623), .A(n272), .ZN(\U27/Z_4 ) );
  OAI21_X2 U560 ( .B1(n1665), .B2(n1623), .A(n266), .ZN(\U28/Z_0 ) );
  OAI21_X2 U561 ( .B1(n49), .B2(n1623), .A(n282), .ZN(\U27/Z_0 ) );
  OAI21_X2 U562 ( .B1(n43), .B2(n1623), .A(n270), .ZN(\U27/Z_6 ) );
  OAI21_X2 U563 ( .B1(n42), .B2(n1365), .A(n269), .ZN(\U27/Z_7 ) );
  OAI21_X2 U564 ( .B1(n1365), .B2(n66), .A(n265), .ZN(\U29/Z_0 ) );
  OAI21_X2 U565 ( .B1(n1365), .B2(n65), .A(n264), .ZN(\U29/Z_1 ) );
  OAI21_X2 U566 ( .B1(n1365), .B2(n64), .A(n257), .ZN(\U29/Z_2 ) );
  OAI21_X2 U567 ( .B1(n1365), .B2(n63), .A(n256), .ZN(\U29/Z_3 ) );
  OAI21_X2 U568 ( .B1(n1365), .B2(n62), .A(n255), .ZN(\U29/Z_4 ) );
  OAI21_X2 U569 ( .B1(n1623), .B2(n61), .A(n254), .ZN(\U29/Z_5 ) );
  OAI21_X2 U570 ( .B1(n1365), .B2(n60), .A(n253), .ZN(\U29/Z_6 ) );
  OAI21_X2 U571 ( .B1(n1623), .B2(n59), .A(n252), .ZN(\U29/Z_7 ) );
  OAI21_X2 U572 ( .B1(n48), .B2(n1365), .A(n281), .ZN(\U27/Z_1 ) );
  OAI21_X2 U573 ( .B1(n46), .B2(n1365), .A(n273), .ZN(\U27/Z_3 ) );
  OAI21_X2 U574 ( .B1(n67), .B2(n1365), .A(n289), .ZN(\U26/Z_35 ) );
  OR2_X1 U575 ( .A1(n1635), .A2(\U14/DATA1_27 ), .ZN(n1469) );
  OR2_X1 U576 ( .A1(n1635), .A2(\U14/DATA1_25 ), .ZN(n1471) );
  BUF_X4 U577 ( .A(inputBaseOffset), .Z(m1ReadAddr[15]) );
  XOR2_X1 U578 ( .A(n1798), .B(n1839), .Z(\U14/DATA1_21 ) );
  OR2_X1 U579 ( .A1(n1619), .A2(n1852), .ZN(n1618) );
  INV_X4 U580 ( .A(n1859), .ZN(n1619) );
  NOR2_X2 U581 ( .A1(n1800), .A2(n1621), .ZN(n1620) );
  XNOR2_X1 U582 ( .A(n1712), .B(\U3/U1/Z_0 ), .ZN(n1676) );
  INV_X2 U583 ( .A(n1862), .ZN(n1864) );
  XNOR2_X1 U584 ( .A(\U27/DATA2_1 ), .B(\U29/DATA2_1 ), .ZN(n1653) );
  AND2_X1 U585 ( .A1(\U16/DATA1_0 ), .A2(start), .ZN(\U16/Z_0 ) );
  NOR2_X2 U586 ( .A1(n404), .A2(n1369), .ZN(n1638) );
  AOI221_X2 U587 ( .B1(n337), .B2(\U13/DATA1_3 ), .C1(n339), .C2(n369), .A(
        n1638), .ZN(n362) );
  INV_X4 U588 ( .A(\U15/DATA1_4 ), .ZN(n1664) );
  NOR2_X2 U589 ( .A1(n1635), .A2(n1664), .ZN(\U15/Z_4 ) );
  INV_X4 U590 ( .A(n369), .ZN(n1648) );
  NAND2_X2 U591 ( .A1(n409), .A2(\U13/DATA1_3 ), .ZN(n1639) );
  OAI221_X2 U592 ( .B1(n333), .B2(n1648), .C1(n408), .C2(n1369), .A(n1639), 
        .ZN(n1640) );
  INV_X4 U593 ( .A(\U15/DATA1_5 ), .ZN(n1663) );
  NOR2_X2 U594 ( .A1(n1635), .A2(n1663), .ZN(\U15/Z_5 ) );
  NOR2_X2 U595 ( .A1(n386), .A2(n1369), .ZN(n1641) );
  AOI221_X2 U596 ( .B1(n322), .B2(\U13/DATA1_3 ), .C1(n323), .C2(n369), .A(
        n1641), .ZN(n350) );
  NOR2_X2 U597 ( .A1(n1635), .A2(n1372), .ZN(\U15/Z_6 ) );
  AND2_X1 U598 ( .A1(n435), .A2(n436), .ZN(n344) );
  NOR2_X2 U599 ( .A1(n1635), .A2(n1373), .ZN(\U15/Z_7 ) );
  NOR2_X2 U600 ( .A1(n371), .A2(n1369), .ZN(n1642) );
  AOI221_X2 U601 ( .B1(n351), .B2(n369), .C1(n352), .C2(\U13/DATA1_3 ), .A(
        n1642), .ZN(n368) );
  INV_X4 U602 ( .A(\U15/DATA1_2 ), .ZN(n1666) );
  NOR2_X2 U603 ( .A1(n1635), .A2(n1666), .ZN(\U15/Z_2 ) );
  NOR2_X2 U604 ( .A1(n427), .A2(n1369), .ZN(n1643) );
  AOI221_X2 U605 ( .B1(n346), .B2(n369), .C1(n345), .C2(\U13/DATA1_3 ), .A(
        n1643), .ZN(n426) );
  INV_X4 U606 ( .A(\U15/DATA1_3 ), .ZN(n1667) );
  NOR2_X2 U607 ( .A1(n1635), .A2(n1667), .ZN(\U15/Z_3 ) );
  NAND2_X2 U608 ( .A1(n393), .A2(\U13/DATA1_3 ), .ZN(n1644) );
  OAI221_X2 U609 ( .B1(n365), .B2(n1648), .C1(n389), .C2(n1369), .A(n1644), 
        .ZN(n1645) );
  NOR2_X2 U610 ( .A1(n1635), .A2(n1646), .ZN(\U15/Z_0 ) );
  NAND2_X2 U611 ( .A1(n418), .A2(\U13/DATA1_3 ), .ZN(n1647) );
  OAI221_X2 U612 ( .B1(n359), .B2(n1648), .C1(n417), .C2(n1369), .A(n1647), 
        .ZN(n1649) );
  NOR2_X2 U613 ( .A1(n1635), .A2(n1374), .ZN(\U15/Z_1 ) );
  INV_X4 U614 ( .A(\U25/DATA2_0 ), .ZN(n1662) );
  XNOR2_X2 U615 ( .A(n61), .B(\U27/DATA2_5 ), .ZN(n1651) );
  XNOR2_X2 U616 ( .A(n62), .B(\U27/DATA2_4 ), .ZN(n1650) );
  NOR3_X2 U617 ( .A1(n1665), .A2(n1651), .A3(n1650), .ZN(n1661) );
  XNOR2_X2 U618 ( .A(\U27/DATA2_0 ), .B(\U29/DATA2_0 ), .ZN(n1652) );
  NAND2_X2 U619 ( .A1(n1653), .A2(n1652), .ZN(n1656) );
  XNOR2_X2 U620 ( .A(n64), .B(\U27/DATA2_2 ), .ZN(n1655) );
  XNOR2_X2 U621 ( .A(n63), .B(\U27/DATA2_3 ), .ZN(n1654) );
  NOR3_X2 U622 ( .A1(n1656), .A2(n1655), .A3(n1654), .ZN(n1660) );
  XNOR2_X2 U623 ( .A(\U27/DATA2_6 ), .B(n60), .ZN(n1658) );
  XNOR2_X2 U624 ( .A(\U27/DATA2_7 ), .B(n59), .ZN(n1657) );
  NOR2_X2 U625 ( .A1(n1658), .A2(n1657), .ZN(n1659) );
  OAI22_X2 U626 ( .A1(n1772), .A2(n1662), .B1(n102), .B2(n1627), .ZN(\U18/Z_0 ) );
  XOR2_X2 U627 ( .A(n42), .B(\U15/DATA1_7 ), .Z(n1671) );
  XOR2_X2 U628 ( .A(n43), .B(\U15/DATA1_6 ), .Z(n1670) );
  NAND2_X2 U629 ( .A1(n1631), .A2(n1673), .ZN(n1674) );
  NAND2_X2 U630 ( .A1(n318), .A2(n1674), .ZN(\U26/Z_0 ) );
  INV_X4 U631 ( .A(\U25/DATA2_1 ), .ZN(n1675) );
  OAI22_X2 U632 ( .A1(n1772), .A2(n1675), .B1(n101), .B2(n1627), .ZN(\U18/Z_1 ) );
  MUX2_X2 U633 ( .A(\U3/U1/DATA1_1 ), .B(n1677), .S(n1871), .Z(n1712) );
  NOR2_X2 U634 ( .A1(n1635), .A2(n1676), .ZN(\U14/Z_1 ) );
  NAND2_X2 U635 ( .A1(n1631), .A2(n1677), .ZN(n1678) );
  NAND2_X2 U636 ( .A1(n317), .A2(n1678), .ZN(\U26/Z_1 ) );
  INV_X4 U637 ( .A(\U25/DATA2_2 ), .ZN(n1679) );
  OAI22_X2 U638 ( .A1(n1772), .A2(n1679), .B1(n100), .B2(n1627), .ZN(\U18/Z_2 ) );
  MUX2_X2 U639 ( .A(\U3/U1/DATA1_2 ), .B(n1681), .S(n1871), .Z(n1684) );
  INV_X4 U640 ( .A(n1684), .ZN(n1716) );
  XOR2_X2 U641 ( .A(n1716), .B(n1451), .Z(n1680) );
  NOR2_X2 U642 ( .A1(n1635), .A2(n1680), .ZN(\U14/Z_2 ) );
  NAND2_X2 U643 ( .A1(n1631), .A2(n1681), .ZN(n1682) );
  NAND2_X2 U644 ( .A1(n306), .A2(n1682), .ZN(\U26/Z_2 ) );
  INV_X4 U645 ( .A(\U25/DATA2_3 ), .ZN(n1683) );
  OAI22_X2 U646 ( .A1(n1772), .A2(n1683), .B1(n99), .B2(n1627), .ZN(\U18/Z_3 )
         );
  MUX2_X2 U647 ( .A(\U3/U1/DATA1_3 ), .B(n1686), .S(n1871), .Z(n1713) );
  NOR2_X2 U648 ( .A1(n1635), .A2(n1685), .ZN(\U14/Z_3 ) );
  NAND2_X2 U649 ( .A1(n1631), .A2(n1686), .ZN(n1687) );
  NAND2_X2 U650 ( .A1(n295), .A2(n1687), .ZN(\U26/Z_3 ) );
  INV_X4 U651 ( .A(\U25/DATA2_4 ), .ZN(n1688) );
  OAI22_X2 U652 ( .A1(n1772), .A2(n1688), .B1(n98), .B2(n1627), .ZN(\U18/Z_4 )
         );
  MUX2_X2 U653 ( .A(\U3/U1/DATA1_4 ), .B(n1690), .S(n1871), .Z(n1693) );
  INV_X4 U654 ( .A(n1693), .ZN(n1715) );
  XOR2_X2 U655 ( .A(n1715), .B(n1461), .Z(n1689) );
  NOR2_X2 U656 ( .A1(n1635), .A2(n1689), .ZN(\U14/Z_4 ) );
  NAND2_X2 U657 ( .A1(n1631), .A2(n1690), .ZN(n1691) );
  NAND2_X2 U658 ( .A1(n288), .A2(n1691), .ZN(\U26/Z_4 ) );
  INV_X4 U659 ( .A(\U25/DATA2_5 ), .ZN(n1692) );
  OAI22_X2 U660 ( .A1(n1772), .A2(n1692), .B1(n97), .B2(n1627), .ZN(\U18/Z_5 )
         );
  MUX2_X2 U661 ( .A(\U3/U1/DATA1_5 ), .B(n1695), .S(n1871), .Z(n1714) );
  XNOR2_X2 U662 ( .A(n1714), .B(n1459), .ZN(n1694) );
  NOR2_X2 U663 ( .A1(n1635), .A2(n1694), .ZN(\U14/Z_5 ) );
  NAND2_X2 U664 ( .A1(n1631), .A2(n1695), .ZN(n1696) );
  NAND2_X2 U665 ( .A1(n287), .A2(n1696), .ZN(\U26/Z_5 ) );
  INV_X4 U666 ( .A(\U25/DATA2_6 ), .ZN(n1697) );
  OAI22_X2 U667 ( .A1(n1772), .A2(n1697), .B1(n96), .B2(n1627), .ZN(\U18/Z_6 )
         );
  MUX2_X2 U668 ( .A(\U3/U1/DATA1_6 ), .B(n1699), .S(n1871), .Z(n1718) );
  XNOR2_X2 U669 ( .A(n1718), .B(n1455), .ZN(n1698) );
  NOR2_X2 U670 ( .A1(n1635), .A2(n1698), .ZN(\U14/Z_6 ) );
  NAND2_X2 U671 ( .A1(n1631), .A2(n1699), .ZN(n1700) );
  NAND2_X2 U672 ( .A1(n286), .A2(n1700), .ZN(\U26/Z_6 ) );
  INV_X4 U673 ( .A(\U25/DATA2_7 ), .ZN(n1701) );
  OAI22_X2 U674 ( .A1(n1772), .A2(n1701), .B1(n95), .B2(n1627), .ZN(\U18/Z_7 )
         );
  MUX2_X2 U675 ( .A(\U3/U1/DATA1_7 ), .B(n1703), .S(n1871), .Z(n1719) );
  NAND2_X2 U676 ( .A1(n1455), .A2(n1718), .ZN(n1706) );
  XNOR2_X2 U677 ( .A(n1443), .B(n1706), .ZN(n1702) );
  NOR2_X2 U678 ( .A1(n1635), .A2(n1702), .ZN(\U14/Z_7 ) );
  NAND2_X2 U679 ( .A1(n1631), .A2(n1703), .ZN(n1704) );
  NAND2_X2 U680 ( .A1(n285), .A2(n1704), .ZN(\U26/Z_7 ) );
  INV_X4 U681 ( .A(\U25/DATA2_8 ), .ZN(n1705) );
  OAI22_X2 U682 ( .A1(n1772), .A2(n1705), .B1(n94), .B2(n1627), .ZN(\U18/Z_8 )
         );
  MUX2_X2 U683 ( .A(\U3/U1/DATA1_8 ), .B(n1709), .S(n1871), .Z(n1717) );
  NOR2_X2 U684 ( .A1(n1443), .A2(n1706), .ZN(n1707) );
  NOR2_X2 U685 ( .A1(n1635), .A2(n1708), .ZN(\U14/Z_8 ) );
  NAND2_X2 U686 ( .A1(n1631), .A2(n1709), .ZN(n1710) );
  NAND2_X2 U687 ( .A1(n284), .A2(n1710), .ZN(\U26/Z_8 ) );
  INV_X4 U688 ( .A(\U25/DATA2_9 ), .ZN(n1711) );
  OAI22_X2 U689 ( .A1(n1772), .A2(n1711), .B1(n93), .B2(n1627), .ZN(\U18/Z_9 )
         );
  MUX2_X2 U690 ( .A(\U3/U1/DATA1_9 ), .B(n1721), .S(n1871), .Z(n1747) );
  NOR2_X2 U691 ( .A1(n1635), .A2(n1720), .ZN(\U14/Z_9 ) );
  NAND2_X2 U692 ( .A1(n1631), .A2(n1721), .ZN(n1722) );
  NAND2_X2 U693 ( .A1(n283), .A2(n1722), .ZN(\U26/Z_9 ) );
  INV_X4 U694 ( .A(\U25/DATA2_10 ), .ZN(n1723) );
  OAI22_X2 U695 ( .A1(n1772), .A2(n1723), .B1(n92), .B2(n1627), .ZN(\U18/Z_10 ) );
  MUX2_X2 U696 ( .A(\U3/U1/DATA1_10 ), .B(n1725), .S(n1871), .Z(n1751) );
  XNOR2_X2 U697 ( .A(n1751), .B(n1456), .ZN(n1724) );
  NOR2_X2 U698 ( .A1(n1635), .A2(n1724), .ZN(\U14/Z_10 ) );
  NAND2_X2 U704 ( .A1(n1631), .A2(n1725), .ZN(n1726) );
  NAND2_X2 U707 ( .A1(n316), .A2(n1726), .ZN(\U26/Z_10 ) );
  INV_X4 U709 ( .A(\U25/DATA2_11 ), .ZN(n1727) );
  OAI22_X2 U710 ( .A1(n1772), .A2(n1727), .B1(n91), .B2(n1627), .ZN(\U18/Z_11 ) );
  MUX2_X2 U711 ( .A(\U3/U1/DATA1_11 ), .B(n1729), .S(n1871), .Z(n1752) );
  XNOR2_X2 U712 ( .A(n1752), .B(n1452), .ZN(n1728) );
  NOR2_X2 U713 ( .A1(n1635), .A2(n1728), .ZN(\U14/Z_11 ) );
  NAND2_X2 U714 ( .A1(n1631), .A2(n1729), .ZN(n1730) );
  NAND2_X2 U715 ( .A1(n315), .A2(n1730), .ZN(\U26/Z_11 ) );
  INV_X4 U716 ( .A(\U25/DATA2_12 ), .ZN(n1731) );
  OAI22_X2 U717 ( .A1(n1772), .A2(n1731), .B1(n90), .B2(n1627), .ZN(\U18/Z_12 ) );
  MUX2_X2 U718 ( .A(\U3/U1/DATA1_12 ), .B(n1733), .S(n1629), .Z(n1753) );
  XNOR2_X2 U719 ( .A(n1753), .B(n1454), .ZN(n1732) );
  NOR2_X2 U720 ( .A1(n1635), .A2(n1732), .ZN(\U14/Z_12 ) );
  NAND2_X2 U721 ( .A1(n1631), .A2(n1733), .ZN(n1734) );
  NAND2_X2 U722 ( .A1(n314), .A2(n1734), .ZN(\U26/Z_12 ) );
  INV_X4 U723 ( .A(\U25/DATA2_13 ), .ZN(n1735) );
  OAI22_X2 U724 ( .A1(n1772), .A2(n1735), .B1(n89), .B2(n1627), .ZN(\U18/Z_13 ) );
  MUX2_X2 U725 ( .A(\U3/U1/DATA1_13 ), .B(n1737), .S(n1871), .Z(n1748) );
  INV_X4 U726 ( .A(n1748), .ZN(n1741) );
  NAND2_X2 U727 ( .A1(n1454), .A2(n1753), .ZN(n1740) );
  XNOR2_X2 U728 ( .A(n1741), .B(n1740), .ZN(n1736) );
  NOR2_X2 U729 ( .A1(n1635), .A2(n1736), .ZN(\U14/Z_13 ) );
  NAND2_X2 U730 ( .A1(n1631), .A2(n1737), .ZN(n1738) );
  NAND2_X2 U731 ( .A1(n313), .A2(n1738), .ZN(\U26/Z_13 ) );
  INV_X4 U732 ( .A(\U25/DATA2_14 ), .ZN(n1739) );
  OAI22_X2 U733 ( .A1(n1772), .A2(n1739), .B1(n88), .B2(n1627), .ZN(\U18/Z_14 ) );
  MUX2_X2 U734 ( .A(\U3/U1/DATA1_14 ), .B(n1744), .S(n1871), .Z(n1749) );
  NOR2_X2 U735 ( .A1(n1741), .A2(n1740), .ZN(n1742) );
  NOR2_X2 U736 ( .A1(n1635), .A2(n1743), .ZN(\U14/Z_14 ) );
  NAND2_X2 U737 ( .A1(n1631), .A2(n1744), .ZN(n1745) );
  NAND2_X2 U738 ( .A1(n312), .A2(n1745), .ZN(\U26/Z_14 ) );
  INV_X4 U739 ( .A(\U25/DATA2_15 ), .ZN(n1746) );
  OAI22_X2 U740 ( .A1(n1772), .A2(n1746), .B1(n87), .B2(n1627), .ZN(\U18/Z_15 ) );
  MUX2_X2 U741 ( .A(\U3/U1/DATA1_15 ), .B(n1756), .S(n1628), .Z(n1788) );
  NAND3_X2 U742 ( .A1(n1749), .A2(n1748), .A3(n1747), .ZN(n1750) );
  INV_X4 U743 ( .A(n1750), .ZN(n1782) );
  INV_X4 U744 ( .A(n1785), .ZN(n1754) );
  XNOR2_X2 U745 ( .A(n1788), .B(n1448), .ZN(n1755) );
  NOR2_X2 U746 ( .A1(n1635), .A2(n1755), .ZN(\U14/Z_15 ) );
  NAND2_X2 U747 ( .A1(n1631), .A2(n1756), .ZN(n1757) );
  NAND2_X2 U748 ( .A1(n311), .A2(n1757), .ZN(\U26/Z_15 ) );
  INV_X4 U749 ( .A(\U25/DATA2_16 ), .ZN(n1758) );
  OAI22_X2 U750 ( .A1(n1772), .A2(n1758), .B1(n86), .B2(n1627), .ZN(\U18/Z_16 ) );
  MUX2_X2 U751 ( .A(\U3/U1/DATA1_16 ), .B(n1760), .S(n1628), .Z(n1763) );
  INV_X4 U752 ( .A(n1763), .ZN(n1783) );
  XOR2_X2 U753 ( .A(n1783), .B(n1460), .Z(n1759) );
  NOR2_X2 U754 ( .A1(n1635), .A2(n1759), .ZN(\U14/Z_16 ) );
  NAND2_X2 U755 ( .A1(n1631), .A2(n1760), .ZN(n1761) );
  NAND2_X2 U756 ( .A1(n310), .A2(n1761), .ZN(\U26/Z_16 ) );
  INV_X4 U757 ( .A(\U25/DATA2_17 ), .ZN(n1762) );
  OAI22_X2 U758 ( .A1(n1772), .A2(n1762), .B1(n85), .B2(n1627), .ZN(\U18/Z_17 ) );
  MUX2_X2 U759 ( .A(\U3/U1/DATA1_17 ), .B(n1765), .S(n1629), .Z(n1781) );
  NOR2_X2 U760 ( .A1(n1635), .A2(n1764), .ZN(\U14/Z_17 ) );
  NAND2_X2 U761 ( .A1(n1631), .A2(n1765), .ZN(n1766) );
  NAND2_X2 U762 ( .A1(n309), .A2(n1766), .ZN(\U26/Z_17 ) );
  INV_X4 U763 ( .A(\U25/DATA2_18 ), .ZN(n1767) );
  OAI22_X2 U764 ( .A1(n1772), .A2(n1767), .B1(n84), .B2(n1627), .ZN(\U18/Z_18 ) );
  MUX2_X2 U765 ( .A(\U3/U1/DATA1_18 ), .B(n1769), .S(n1629), .Z(n1794) );
  XNOR2_X2 U766 ( .A(n1794), .B(n1453), .ZN(n1768) );
  NOR2_X2 U767 ( .A1(n1635), .A2(n1768), .ZN(\U14/Z_18 ) );
  NAND2_X2 U768 ( .A1(n1631), .A2(n1769), .ZN(n1770) );
  NAND2_X2 U769 ( .A1(n308), .A2(n1770), .ZN(\U26/Z_18 ) );
  INV_X4 U770 ( .A(\U25/DATA2_19 ), .ZN(n1771) );
  OAI22_X2 U771 ( .A1(n1772), .A2(n1771), .B1(n83), .B2(n1627), .ZN(\U18/Z_19 ) );
  MUX2_X2 U772 ( .A(\U3/U1/DATA1_19 ), .B(n1775), .S(n1628), .Z(n1773) );
  INV_X4 U773 ( .A(n1773), .ZN(n1786) );
  NOR2_X2 U774 ( .A1(n1635), .A2(n1774), .ZN(\U14/Z_19 ) );
  NAND2_X2 U775 ( .A1(n1631), .A2(n1775), .ZN(n1776) );
  NAND2_X2 U776 ( .A1(n307), .A2(n1776), .ZN(\U26/Z_19 ) );
  NOR2_X2 U777 ( .A1(n82), .A2(n1627), .ZN(\U18/Z_20 ) );
  MUX2_X2 U778 ( .A(\U3/U1/DATA1_20 ), .B(n1779), .S(n1628), .Z(n1789) );
  NAND2_X2 U779 ( .A1(n1631), .A2(n1779), .ZN(n1780) );
  NAND2_X2 U780 ( .A1(n305), .A2(n1780), .ZN(\U26/Z_20 ) );
  NAND2_X2 U781 ( .A1(n81), .A2(n1360), .ZN(\U18/Z_21 ) );
  INV_X4 U782 ( .A(n1788), .ZN(n1791) );
  INV_X4 U783 ( .A(n1789), .ZN(n1790) );
  NOR2_X2 U784 ( .A1(n1791), .A2(n1790), .ZN(n1792) );
  MUX2_X2 U785 ( .A(\U3/U1/DATA1_21 ), .B(n1796), .S(n1629), .Z(n1799) );
  INV_X4 U786 ( .A(n1799), .ZN(n1839) );
  NAND2_X2 U787 ( .A1(n1631), .A2(n1796), .ZN(n1797) );
  NAND2_X2 U788 ( .A1(n304), .A2(n1797), .ZN(\U26/Z_21 ) );
  NOR2_X2 U789 ( .A1(n80), .A2(n1627), .ZN(\U18/Z_22 ) );
  MUX2_X2 U790 ( .A(\U3/U1/DATA1_22 ), .B(n1802), .S(n1871), .Z(n1834) );
  INV_X4 U791 ( .A(n1439), .ZN(n1842) );
  NAND2_X2 U792 ( .A1(n1842), .A2(n1799), .ZN(n1800) );
  NOR2_X2 U793 ( .A1(n1635), .A2(n1801), .ZN(\U14/Z_22 ) );
  NAND2_X2 U794 ( .A1(n1631), .A2(n1802), .ZN(n1803) );
  NAND2_X2 U795 ( .A1(n303), .A2(n1803), .ZN(\U26/Z_22 ) );
  NAND2_X2 U796 ( .A1(n79), .A2(n1360), .ZN(\U18/Z_23 ) );
  MUX2_X2 U797 ( .A(\U3/U1/DATA1_23 ), .B(n1804), .S(n1628), .Z(n1806) );
  INV_X4 U798 ( .A(n1806), .ZN(n1838) );
  NAND2_X2 U799 ( .A1(n1631), .A2(n1804), .ZN(n1805) );
  NAND2_X2 U800 ( .A1(n302), .A2(n1805), .ZN(\U26/Z_23 ) );
  NOR2_X2 U801 ( .A1(n78), .A2(n1627), .ZN(\U18/Z_24 ) );
  MUX2_X2 U802 ( .A(\U3/U1/DATA1_24 ), .B(n1808), .S(n1628), .Z(n1835) );
  INV_X4 U803 ( .A(n1824), .ZN(n1810) );
  XNOR2_X2 U804 ( .A(n1835), .B(n1810), .ZN(n1807) );
  NOR2_X2 U805 ( .A1(n1635), .A2(n1807), .ZN(\U14/Z_24 ) );
  NAND2_X2 U806 ( .A1(n1631), .A2(n1808), .ZN(n1809) );
  NAND2_X2 U807 ( .A1(n301), .A2(n1809), .ZN(\U26/Z_24 ) );
  NAND2_X2 U808 ( .A1(n77), .A2(n1360), .ZN(\U18/Z_25 ) );
  NAND2_X2 U809 ( .A1(n1810), .A2(n1835), .ZN(n1813) );
  MUX2_X2 U810 ( .A(\U3/U1/DATA1_25 ), .B(n1811), .S(n1628), .Z(n1819) );
  NAND2_X2 U811 ( .A1(n1633), .A2(n1811), .ZN(n1812) );
  NAND2_X2 U812 ( .A1(n300), .A2(n1812), .ZN(\U26/Z_25 ) );
  NOR2_X2 U813 ( .A1(n76), .A2(n1627), .ZN(\U18/Z_26 ) );
  MUX2_X2 U814 ( .A(\U3/U1/DATA1_26 ), .B(n1816), .S(n1628), .Z(n1836) );
  INV_X4 U815 ( .A(n1836), .ZN(n1828) );
  INV_X4 U816 ( .A(n1813), .ZN(n1814) );
  XNOR2_X2 U817 ( .A(n1828), .B(n1827), .ZN(n1815) );
  NOR2_X2 U818 ( .A1(n1635), .A2(n1815), .ZN(\U14/Z_26 ) );
  NAND2_X2 U819 ( .A1(n1633), .A2(n1816), .ZN(n1817) );
  NAND2_X2 U820 ( .A1(n299), .A2(n1817), .ZN(\U26/Z_26 ) );
  NAND2_X2 U821 ( .A1(n75), .A2(n1360), .ZN(\U18/Z_27 ) );
  MUX2_X2 U822 ( .A(\U3/U1/DATA1_27 ), .B(n1825), .S(n1871), .Z(n1820) );
  INV_X4 U823 ( .A(n1820), .ZN(n1829) );
  NAND2_X2 U824 ( .A1(n1835), .A2(n1836), .ZN(n1821) );
  INV_X4 U825 ( .A(n1821), .ZN(n1818) );
  NAND2_X2 U826 ( .A1(n1818), .A2(n1819), .ZN(n1823) );
  NAND2_X2 U827 ( .A1(n1820), .A2(n1819), .ZN(n1840) );
  NOR3_X2 U828 ( .A1(n1824), .A2(n1840), .A3(n1821), .ZN(n1822) );
  AOI221_X2 U829 ( .B1(n1829), .B2(n1824), .C1(n1829), .C2(n1823), .A(n1822), 
        .ZN(\U14/DATA1_27 ) );
  NAND2_X2 U830 ( .A1(n1633), .A2(n1825), .ZN(n1826) );
  NAND2_X2 U831 ( .A1(n298), .A2(n1826), .ZN(\U26/Z_27 ) );
  NOR2_X2 U832 ( .A1(n74), .A2(n1627), .ZN(\U18/Z_28 ) );
  MUX2_X2 U833 ( .A(\U3/U1/DATA1_28 ), .B(n1832), .S(n1628), .Z(n1837) );
  NOR2_X2 U834 ( .A1(n1635), .A2(n1831), .ZN(\U14/Z_28 ) );
  NAND2_X2 U835 ( .A1(n1633), .A2(n1832), .ZN(n1833) );
  NAND2_X2 U836 ( .A1(n297), .A2(n1833), .ZN(\U26/Z_28 ) );
  NAND2_X2 U837 ( .A1(n73), .A2(n1360), .ZN(\U18/Z_29 ) );
  NAND4_X2 U838 ( .A1(n1837), .A2(n1836), .A3(n1835), .A4(n1834), .ZN(n1841)
         );
  NOR4_X2 U839 ( .A1(n1841), .A2(n1840), .A3(n1839), .A4(n1838), .ZN(n1843) );
  NAND2_X2 U840 ( .A1(n1843), .A2(n1842), .ZN(n1846) );
  MUX2_X2 U841 ( .A(\U3/U1/DATA1_29 ), .B(n1844), .S(n1628), .Z(n1847) );
  NAND2_X2 U842 ( .A1(n1633), .A2(n1844), .ZN(n1845) );
  NAND2_X2 U843 ( .A1(n296), .A2(n1845), .ZN(\U26/Z_29 ) );
  NOR2_X2 U844 ( .A1(n72), .A2(n1627), .ZN(\U18/Z_30 ) );
  MUX2_X2 U845 ( .A(\U3/U1/DATA1_30 ), .B(n1849), .S(n1628), .Z(n1851) );
  NOR2_X2 U846 ( .A1(n1635), .A2(n1848), .ZN(\U14/Z_30 ) );
  NAND2_X2 U847 ( .A1(n1633), .A2(n1849), .ZN(n1850) );
  NAND2_X2 U848 ( .A1(n294), .A2(n1850), .ZN(\U26/Z_30 ) );
  NAND2_X2 U849 ( .A1(n71), .A2(n1360), .ZN(\U18/Z_31 ) );
  MUX2_X2 U850 ( .A(\U3/U1/DATA1_31 ), .B(n1364), .S(n1629), .Z(n1855) );
  INV_X4 U851 ( .A(n1855), .ZN(n1852) );
  NAND2_X2 U852 ( .A1(n1633), .A2(n1364), .ZN(n1853) );
  NAND2_X2 U853 ( .A1(n293), .A2(n1853), .ZN(\U26/Z_31 ) );
  NOR2_X2 U854 ( .A1(n70), .A2(n1627), .ZN(\U18/Z_32 ) );
  MUX2_X2 U855 ( .A(\U3/U1/DATA1_32 ), .B(n1857), .S(n1629), .Z(n1859) );
  XNOR2_X2 U856 ( .A(n1859), .B(n1622), .ZN(n1856) );
  NOR2_X2 U857 ( .A1(n1635), .A2(n1856), .ZN(\U14/Z_32 ) );
  NAND2_X2 U858 ( .A1(n1631), .A2(n1857), .ZN(n1858) );
  NAND2_X2 U859 ( .A1(n292), .A2(n1858), .ZN(\U26/Z_32 ) );
  NAND2_X2 U860 ( .A1(n69), .A2(n1360), .ZN(\U18/Z_33 ) );
  MUX2_X2 U861 ( .A(\U3/U1/DATA1_33 ), .B(n1860), .S(n1629), .Z(n1863) );
  NAND2_X2 U862 ( .A1(n1631), .A2(n1860), .ZN(n1861) );
  NAND2_X2 U863 ( .A1(n291), .A2(n1861), .ZN(\U26/Z_33 ) );
  NOR2_X2 U864 ( .A1(n68), .A2(n1627), .ZN(\U18/Z_34 ) );
  MUX2_X2 U865 ( .A(\U3/U1/DATA1_34 ), .B(n1867), .S(n1629), .Z(n1869) );
  NAND2_X2 U866 ( .A1(n1864), .A2(n1863), .ZN(n1865) );
  INV_X4 U867 ( .A(n1865), .ZN(n1870) );
  XNOR2_X2 U868 ( .A(n1869), .B(n1870), .ZN(n1866) );
  NOR2_X2 U869 ( .A1(n1635), .A2(n1866), .ZN(\U14/Z_34 ) );
  NAND2_X2 U870 ( .A1(n1631), .A2(n1867), .ZN(n1868) );
  NAND2_X2 U871 ( .A1(n290), .A2(n1868), .ZN(\U26/Z_34 ) );
  NAND2_X2 U872 ( .A1(n67), .A2(n1360), .ZN(\U18/Z_35 ) );
  NAND2_X2 U873 ( .A1(n1870), .A2(n1869), .ZN(n1873) );
  MUX2_X2 U874 ( .A(\U3/U1/DATA1_35 ), .B(\U3/U1/DATA2_35 ), .S(n1628), .Z(
        n1872) );
  NAND2_X2 U875 ( .A1(n1634), .A2(n1874), .ZN(\U14/Z_35 ) );
  NAND2_X2 U876 ( .A1(n340), .A2(n1359), .ZN(n1882) );
  INV_X4 U877 ( .A(n1882), .ZN(n1875) );
  NAND3_X2 U878 ( .A1(\U5/DATA1_1 ), .A2(\U5/DATA1_0 ), .A3(\U5/DATA1_2 ), 
        .ZN(n1890) );
  INV_X4 U879 ( .A(n1890), .ZN(n1893) );
  NAND3_X2 U880 ( .A1(\U5/DATA1_4 ), .A2(\U5/DATA1_3 ), .A3(n1893), .ZN(n1899)
         );
  INV_X4 U881 ( .A(n1899), .ZN(n1902) );
  NAND3_X2 U882 ( .A1(\U5/DATA1_6 ), .A2(\U5/DATA1_5 ), .A3(n1902), .ZN(n1908)
         );
  INV_X4 U883 ( .A(n1908), .ZN(n1916) );
  NOR3_X2 U884 ( .A1(n1878), .A2(n1877), .A3(n1876), .ZN(n1880) );
  NOR4_X2 U885 ( .A1(\U5/DATA1_10 ), .A2(\U5/DATA1_8 ), .A3(\U5/DATA1_13 ), 
        .A4(\U5/DATA1_12 ), .ZN(n1879) );
  NAND4_X2 U886 ( .A1(\U5/DATA1_14 ), .A2(n1916), .A3(n1880), .A4(n1879), .ZN(
        n211) );
  NOR2_X2 U887 ( .A1(n209), .A2(n172), .ZN(n1884) );
  INV_X4 U888 ( .A(n211), .ZN(n1881) );
  NAND2_X2 U889 ( .A1(n1368), .A2(n1881), .ZN(n1883) );
  NAND2_X2 U890 ( .A1(n1882), .A2(n1634), .ZN(n212) );
  INV_X4 U891 ( .A(n209), .ZN(n1926) );
  NAND2_X2 U892 ( .A1(n1926), .A2(n172), .ZN(n1942) );
  NAND2_X2 U893 ( .A1(n1363), .A2(n1942), .ZN(n1886) );
  MUX2_X2 U894 ( .A(n1884), .B(n1886), .S(\U5/DATA1_1 ), .Z(n1943) );
  NAND2_X2 U895 ( .A1(\U5/DATA1_0 ), .A2(n1887), .ZN(n1885) );
  MUX2_X2 U896 ( .A(n1887), .B(n1885), .S(\U5/DATA1_1 ), .Z(n1889) );
  INV_X4 U897 ( .A(n1886), .ZN(n1888) );
  OAI22_X2 U898 ( .A1(n209), .A2(n1889), .B1(n1888), .B2(n1887), .ZN(n1944) );
  NOR2_X2 U899 ( .A1(n209), .A2(n1890), .ZN(n1892) );
  NAND2_X2 U900 ( .A1(n1890), .A2(n1926), .ZN(n1891) );
  NAND2_X2 U901 ( .A1(n1363), .A2(n1891), .ZN(n1895) );
  MUX2_X2 U902 ( .A(n1892), .B(n1895), .S(\U5/DATA1_3 ), .Z(n1945) );
  NAND2_X2 U903 ( .A1(n1893), .A2(n1896), .ZN(n1894) );
  MUX2_X2 U904 ( .A(n1896), .B(n1894), .S(\U5/DATA1_3 ), .Z(n1898) );
  INV_X4 U905 ( .A(n1895), .ZN(n1897) );
  OAI22_X2 U906 ( .A1(n209), .A2(n1898), .B1(n1897), .B2(n1896), .ZN(n1946) );
  NOR2_X2 U907 ( .A1(n209), .A2(n1899), .ZN(n1901) );
  NAND2_X2 U908 ( .A1(n1899), .A2(n1926), .ZN(n1900) );
  NAND2_X2 U909 ( .A1(n1363), .A2(n1900), .ZN(n1904) );
  MUX2_X2 U910 ( .A(n1901), .B(n1904), .S(\U5/DATA1_5 ), .Z(n1947) );
  NAND2_X2 U911 ( .A1(n1902), .A2(n1905), .ZN(n1903) );
  MUX2_X2 U912 ( .A(n1905), .B(n1903), .S(\U5/DATA1_5 ), .Z(n1907) );
  INV_X4 U913 ( .A(n1904), .ZN(n1906) );
  OAI22_X2 U914 ( .A1(n209), .A2(n1907), .B1(n1906), .B2(n1905), .ZN(n1948) );
  NOR2_X2 U915 ( .A1(n209), .A2(n1908), .ZN(n1910) );
  NAND2_X2 U916 ( .A1(n1908), .A2(n1926), .ZN(n1909) );
  NAND2_X2 U917 ( .A1(n1363), .A2(n1909), .ZN(n1912) );
  MUX2_X2 U918 ( .A(n1910), .B(n1912), .S(\U5/DATA1_7 ), .Z(n1949) );
  NAND2_X2 U919 ( .A1(n1916), .A2(n1913), .ZN(n1911) );
  MUX2_X2 U920 ( .A(n1913), .B(n1911), .S(\U5/DATA1_7 ), .Z(n1915) );
  INV_X4 U921 ( .A(n1912), .ZN(n1914) );
  OAI22_X2 U922 ( .A1(n209), .A2(n1915), .B1(n1914), .B2(n1913), .ZN(n1950) );
  NAND3_X2 U923 ( .A1(\U5/DATA1_8 ), .A2(\U5/DATA1_7 ), .A3(n1916), .ZN(n1919)
         );
  NOR2_X2 U924 ( .A1(n209), .A2(n1919), .ZN(n1918) );
  NAND2_X2 U925 ( .A1(n1919), .A2(n1926), .ZN(n1917) );
  NAND2_X2 U926 ( .A1(n1363), .A2(n1917), .ZN(n1921) );
  MUX2_X2 U927 ( .A(n1918), .B(n1921), .S(\U5/DATA1_9 ), .Z(n1951) );
  INV_X4 U928 ( .A(n1919), .ZN(n1925) );
  NAND2_X2 U929 ( .A1(n1925), .A2(n1922), .ZN(n1920) );
  MUX2_X2 U930 ( .A(n1922), .B(n1920), .S(\U5/DATA1_9 ), .Z(n1924) );
  INV_X4 U931 ( .A(n1921), .ZN(n1923) );
  OAI22_X2 U932 ( .A1(n209), .A2(n1924), .B1(n1923), .B2(n1922), .ZN(n1952) );
  NAND3_X2 U933 ( .A1(\U5/DATA1_10 ), .A2(\U5/DATA1_9 ), .A3(n1925), .ZN(n1929) );
  NOR2_X2 U934 ( .A1(n209), .A2(n1929), .ZN(n1928) );
  NAND2_X2 U935 ( .A1(n1929), .A2(n1926), .ZN(n1927) );
  NAND2_X2 U936 ( .A1(n1363), .A2(n1927), .ZN(n1931) );
  MUX2_X2 U937 ( .A(n1928), .B(n1931), .S(\U5/DATA1_11 ), .Z(n1953) );
  INV_X4 U938 ( .A(n1929), .ZN(n1935) );
  NAND2_X2 U939 ( .A1(n1935), .A2(n1932), .ZN(n1930) );
  MUX2_X2 U940 ( .A(n1932), .B(n1930), .S(\U5/DATA1_11 ), .Z(n1934) );
  INV_X4 U941 ( .A(n1931), .ZN(n1933) );
  OAI22_X2 U942 ( .A1(n209), .A2(n1934), .B1(n1933), .B2(n1932), .ZN(n1954) );
  NAND3_X2 U943 ( .A1(\U5/DATA1_12 ), .A2(\U5/DATA1_11 ), .A3(n1935), .ZN(
        n1937) );
  XOR2_X2 U944 ( .A(n1937), .B(\U5/DATA1_13 ), .Z(n1936) );
  OAI22_X2 U945 ( .A1(n209), .A2(n1936), .B1(n1363), .B2(n1463), .ZN(n1955) );
  NAND2_X2 U946 ( .A1(n1368), .A2(n1939), .ZN(n1938) );
  NAND2_X2 U947 ( .A1(n1363), .A2(n1938), .ZN(n1941) );
  NOR2_X2 U948 ( .A1(n209), .A2(n1939), .ZN(n1940) );
  MUX2_X2 U949 ( .A(n1941), .B(n1940), .S(n171), .Z(n510) );
  INV_X4 U950 ( .A(\U12/Z_0 ), .ZN(n1956) );
  INV_X4 U951 ( .A(n434), .ZN(n1957) );
  INV_X4 U952 ( .A(n433), .ZN(n1958) );
  INV_X4 U953 ( .A(n428), .ZN(n1959) );
  INV_X4 U954 ( .A(n422), .ZN(n1960) );
  INV_X4 U955 ( .A(n421), .ZN(n1961) );
  INV_X4 U956 ( .A(n413), .ZN(n1962) );
  INV_X4 U957 ( .A(n412), .ZN(n1963) );
  INV_X4 U958 ( .A(n401), .ZN(n1964) );
  INV_X4 U959 ( .A(n397), .ZN(n1966) );
  INV_X4 U960 ( .A(n396), .ZN(n1967) );
  INV_X4 U961 ( .A(n390), .ZN(n1968) );
  INV_X4 U962 ( .A(n383), .ZN(n1969) );
  INV_X4 U963 ( .A(n379), .ZN(n1971) );
  INV_X4 U964 ( .A(n378), .ZN(n1972) );
  INV_X4 U965 ( .A(n372), .ZN(n1973) );
  INV_X4 U966 ( .A(n425), .ZN(n1974) );
  INV_X4 U967 ( .A(n416), .ZN(n1975) );
  INV_X4 U968 ( .A(n405), .ZN(n1976) );
  INV_X4 U969 ( .A(n387), .ZN(n1977) );
endmodule


module Top ( clock, reset_n, start, M1_ReadBus1, M1_ReadAddress1, M2_ReadBus1, 
        M2_ReadBus2, M2_ReadAddress1, M2_ReadAddress2, M2_WriteBus, 
        M2_WriteAddress, M2_WriteEnable, M3_ReadBus1, M3_ReadBus2, 
        M3_ReadAddress1, M3_ReadAddress2, M3_WriteBus, M3_WriteAddress, 
        M3_WriteEnable, M4_WriteBus, M4_WriteAddress, M4_WriteEnable );
  input [127:0] M1_ReadBus1;
  output [15:0] M1_ReadAddress1;
  input [127:0] M2_ReadBus1;
  input [127:0] M2_ReadBus2;
  output [15:0] M2_ReadAddress1;
  output [15:0] M2_ReadAddress2;
  output [127:0] M2_WriteBus;
  output [15:0] M2_WriteAddress;
  input [127:0] M3_ReadBus1;
  input [127:0] M3_ReadBus2;
  output [15:0] M3_ReadAddress1;
  output [15:0] M3_ReadAddress2;
  output [127:0] M3_WriteBus;
  output [15:0] M3_WriteAddress;
  output [127:0] M4_WriteBus;
  output [15:0] M4_WriteAddress;
  input clock, reset_n, start;
  output M2_WriteEnable, M3_WriteEnable, M4_WriteEnable;
  wire   input_base_offset, output_base_offset, output_start, input_start,
         output_done, input_done, cdf_valid, n16, n17;
  wire   [19:0] cdf_min;
  wire   [19:0] cdf_min_out;
  wire   [19:0] divisor;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  Output_top dut_output_top ( .clock(clock), .reset_n(n16), .start(
        output_start), .CdfMin(cdf_min_out), .divisor(divisor), .M2SP_ReadBus(
        M2_ReadBus2), .M2SP_ReadAddress({M2_ReadAddress2[15], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, M2_ReadAddress2[7:0]}), .M3SP_ReadBus(
        M3_ReadBus2), .M3SP_ReadAddress(M3_ReadAddress2), .WriteEnable(
        M4_WriteEnable), .Output_MEMBus(M4_WriteBus), .Output_MEMAddress(
        M4_WriteAddress), .done(output_done), .output_base_offset(
        output_base_offset) );
  Controllor dut_Controller ( .clock(clock), .reset_n(n16), .start(start), 
        .output_start(output_start), .input_start(input_start), .input_done(
        input_done), .output_done(output_done), .Cdf_Min(cdf_min), 
        .Cdf_Min_Out(cdf_min_out), .Divisor(divisor), .output_base_offset(
        output_base_offset), .input_base_offset(input_base_offset), 
        .cdf_valid(cdf_valid) );
  input_pipeline dut_Input_Pipeline ( .start(input_start), .clock(clock), 
        .rst_n(n16), .m1ReadBus(M1_ReadBus1), .m2ReadBus(M2_ReadBus1), 
        .inputBaseOffset(input_base_offset), .m1ReadAddr(M1_ReadAddress1), 
        .m2ReadAddr(M2_ReadAddress1), .m2WriteAddr(M2_WriteAddress), 
        .m2WriteBus(M2_WriteBus), .m2WE(M2_WriteEnable), .done(input_done), 
        .cdf_min(cdf_min), .cdf_valid(cdf_valid) );
  INV_X4 U1 ( .A(1'b1), .ZN(M2_ReadAddress2[8]) );
  INV_X4 U3 ( .A(1'b1), .ZN(M2_ReadAddress2[9]) );
  INV_X4 U5 ( .A(1'b1), .ZN(M2_ReadAddress2[10]) );
  INV_X4 U7 ( .A(1'b1), .ZN(M2_ReadAddress2[11]) );
  INV_X4 U9 ( .A(1'b1), .ZN(M2_ReadAddress2[12]) );
  INV_X4 U11 ( .A(1'b1), .ZN(M2_ReadAddress2[13]) );
  INV_X4 U13 ( .A(1'b1), .ZN(M2_ReadAddress2[14]) );
  INV_X4 U15 ( .A(n17), .ZN(n16) );
  INV_X4 U16 ( .A(reset_n), .ZN(n17) );
endmodule



module Top(
  input wire clock,
  input wire reset_n,
  input wire start,
  input wire M1_ReadBus1,
  output wire M1_ReadAddress1,
  input wire M2_ReadBus1,
  input wire M2_ReadBus2,
  output wire M2_ReadAddress1,
  output wire M2_ReadAddress2,
  output wire M2_WriteBus,
  output wire M2_WriteAddress,
  output wire M2_WriteEnable,
  input wire M3_ReadBus1,
  output wire M3_ReadAddress1,
  output wire M3_WriteBus,
  output wire M3_WriteAddress,
  output wire M3_WriteEnable,
  output wire M4_WriteBus,
  output wire M4_WriteAddress,
  output wire M4_WriteEnable
  );


  wire input_base_offset, output_base_offset;
  wire output_start, input_start, cdf_start;
  wire output_done,input_done, cdf_done;
  wire [19:0] cdf_min, cdf_min_out, divisor;
  wire cdf_valid;


  Output_top(
    .clock(clock),
    .reset_n(reset_n),
    .start(output_start),
    .CdfMin(cdf_min_out),
    .divisor(divisor),
    .M2SP_ReadBus(M2_ReadBus2),
    .M2SP_ReadAddress(M2_ReadAddress2),
    .M3SP_ReadBus(M3_ReadBus2),
    .M3SP_ReadAddress(M3_ReadAddress2),
    .WriteEnable(M4_WriteEnable),
    .Output_MEMBus(M4_WriteBus),
    .Output_MEMAddress(M4_WriteAddress),
    .done(output_done),
    .output_base_offset(output_base_offset)
    );



  Cdf_top(
    .clock(clock),
    .reset_n(reset_n),
    .start(cdf_start),
    .SP_ReadBus(M2_ReadBus1),
    .SP_ReadAddress(M2_ReadAddress1),
    .WriteEnable(M2_WriteEnable),
    .Output_MEMBus(M2_WriteBus),
    .Output_MEMAddress(M2_WriteAddress),
    .Cdf_Min(cdf_min),
    .done(cdf_done),
    .input_base_offset(input_base_offset),
    .cdf_valid(cdf_valid)
    );



  Controllor(
    .clock(clock),
    .reset_n(reset_n),
    .start(start),
    .output_start(output_start),
    .cdf_start(cdf_start),
    .input_start(input_start),
    .input_done(input_done),
    .output_done(output_done),
    .cdf_done(cdf_done),
    .Cdf_Min(cdf_min),
    .Cdf_Min_Out(cdf_min_out),
    .Divisor(divisor),
    .input_base_offset(input_base_offset),
    .output_base_offset(output_base_offset),
    .cdf_valid(cdf_valid)
    );

//The below module is the first module in the overall pipeline
//This counts how many times each pixel value occurs
  input_pipeline(
    .start(input_start), 
    .clock(clock), 
    .rst_n(reset_n),
    .m1ReadVal(M1_ReadBus), 
    .m2ReadVal(M2_ReadBus),
    .inputBaseOffset(inputBaseOffset),
    .m1ReadAddr(M1_ReadAddress), 
    .m2ReadAddr(M2_ReadAddress), 
    .m2WriteAddr(M2_WriteAddress), 
    .m2WriteVal(M2_Write_Bus),
    .m2WE(M2_WriteEnable),
    .done(input_done)
  );

endmodule
